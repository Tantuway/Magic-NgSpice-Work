* SPICE3 file created from buffer.ext - technology: scmos



.MODEL nfet NMOS VTO=0.7 KP=110U GAMMA=0.4 LAMBDA=0.04 PHI=0.7
.MODEL pfet PMOS VTO=-0.7 KP=50U GAMMA=0.57 LAMBDA=0.05 PHI=0.8
.option scale=1u

M1000 Inverter_0/OUT OUT vdd vdd pfet w=16 l=2
+  ad=144 pd=50 as=288 ps=100
M1001 Inverter_0/OUT OUT gnd Gnd nfet w=8 l=2
+  ad=72 pd=34 as=144 ps=68
M1002 OUT IN vdd vdd pfet w=16 l=2
+  ad=144 pd=50 as=0 ps=0
M1003 OUT IN gnd Gnd nfet w=8 l=2
+  ad=72 pd=34 as=0 ps=0
C0 IN gnd! 7.4fF
C1 OUT gnd! 11.7fF


v3  Inverter_0/OUT  output dc 0 
v2  gnd gnd! dc 0
v1  vdd gnd dc 5
Vin IN gnd pulse(0 5 0 0.1ns 0.1ns 1ns 2ns)
.tran 0.001ns 35.3ns 35.0ns 


.control
run
plot V(output) V(IN) 
.ENDC
.end


