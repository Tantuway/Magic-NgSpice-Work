magic
tech scmos
timestamp 1569346130
<< nwell >>
rect 29 69 64 70
rect 26 62 64 69
rect 29 40 64 62
<< metal1 >>
rect 26 62 64 69
rect 28 34 43 36
rect 28 31 41 34
rect 3 0 63 10
use NAND  NAND_0
timestamp 1569336977
transform 1 0 9 0 1 36
box -8 -34 21 34
use Inverter  Inverter_0
timestamp 1569345144
transform 1 0 44 0 1 37
box -4 -31 20 31
<< end >>
