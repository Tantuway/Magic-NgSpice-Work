* SPICE3 file created from NAND.ext - technology: scmos

.MODEL nfet NMOS VTO=0.7 KP=110U GAMMA=0.4 LAMBDA=0.04 PHI=0.7
.MODEL pfet PMOS VTO=-0.7 KP=50U GAMMA=0.57 LAMBDA=0.05 PHI=0.8

.option scale=1u

M1000 NAND_AB IN_A vdd vdd pfet w=16 l=2
+  ad=192 pd=56 as=160 ps=84
M1001 NAND_AB IN_B  vdd vdd pfet w=16 l=2
+  ad=0 pd=0 as=0 ps=0
M1002 DS IN_A gnd Gnd nfet w=8 l=2
+  ad=96 pd=40 as=40 ps=26
M1003 NAND_AB IN_B DS Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
C0 NAND_AB gnd! 5.3fF
C1 IN_B gnd! 9.8fF
C2 IN_A gnd! 7.3fF


v3 gnd gnd! dc 0V

VDD  vdd gnd DC 5

v2 IN_A gnd PWL (0 0 2N 0 2.1N 5 4N 5 4.1N 0 6N 0 6.1N 5 8N 5 8.1N 0 10N 0 10.1N 5 12N 5 12.1N 0 14N 0 14.1N 5 16N 5 16.1N 0 ) 
v1 IN_B gnd PWL (0 0 4N 0 4.1N 5 8N 5 8.1N 0 12N 0 12.1N 5 16N 5 16.1N 0)

.tran 0.01ns 20ns 0ns 

.control 
run 
plot  V(NAND_AB)
.endc
.end


.control 
run 
plot  V(IN_A)
.endc
.end


.control 
run 
plot  V(IN_B)
.endc
.end

