* SPICE3 file created from /home/mayank/cad/SHIFT_REG_8BIT.ext - technology: scmos

.option scale=1u

M1000 D_Flip_Flop_5/QBAR REG_OUT7 vdd vdd pfet w=16 l=2
+  ad=192 pd=56 as=6272 ps=3088
M1001 vdd D_Flip_Flop_5/NAND_3/IN_B D_Flip_Flop_5/QBAR vdd pfet w=16 l=2
+  ad=0 pd=0 as=0 ps=0
M1002 D_Flip_Flop_5/NAND_3/DS REG_OUT7 gnd Gnd nfet w=8 l=2
+  ad=96 pd=40 as=1856 ps=1104
M1003 D_Flip_Flop_5/QBAR D_Flip_Flop_5/NAND_3/IN_B D_Flip_Flop_5/NAND_3/DS Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1004 D_Flip_Flop_5/NAND_3/IN_B D_Flip_Flop_5/NAND_2/IN_A vdd vdd pfet w=16 l=2
+  ad=192 pd=56 as=0 ps=0
M1005 vdd D_Flip_Flop_3/CLK D_Flip_Flop_5/NAND_3/IN_B vdd pfet w=16 l=2
+  ad=0 pd=0 as=0 ps=0
M1006 D_Flip_Flop_5/NAND_2/DS D_Flip_Flop_5/NAND_2/IN_A gnd Gnd nfet w=8 l=2
+  ad=96 pd=40 as=0 ps=0
M1007 D_Flip_Flop_5/NAND_3/IN_B D_Flip_Flop_3/CLK D_Flip_Flop_5/NAND_2/DS Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1008 D_Flip_Flop_5/NAND_2/IN_A REG_OUT6 vdd vdd pfet w=16 l=2
+  ad=144 pd=50 as=0 ps=0
M1009 D_Flip_Flop_5/NAND_2/IN_A REG_OUT6 gnd Gnd nfet w=8 l=2
+  ad=72 pd=34 as=0 ps=0
M1010 D_Flip_Flop_5/NAND_1/NAND_AB D_Flip_Flop_5/NAND_1/IN_A vdd vdd pfet w=16 l=2
+  ad=192 pd=56 as=0 ps=0
M1011 vdd D_Flip_Flop_5/QBAR D_Flip_Flop_5/NAND_1/NAND_AB vdd pfet w=16 l=2
+  ad=0 pd=0 as=0 ps=0
M1012 D_Flip_Flop_5/NAND_1/DS D_Flip_Flop_5/NAND_1/IN_A gnd Gnd nfet w=8 l=2
+  ad=96 pd=40 as=0 ps=0
M1013 D_Flip_Flop_5/NAND_1/NAND_AB D_Flip_Flop_5/QBAR D_Flip_Flop_5/NAND_1/DS Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1014 D_Flip_Flop_5/NAND_1/IN_A REG_OUT6 vdd vdd pfet w=16 l=2
+  ad=192 pd=56 as=0 ps=0
M1015 vdd D_Flip_Flop_3/CLK D_Flip_Flop_5/NAND_1/IN_A vdd pfet w=16 l=2
+  ad=0 pd=0 as=0 ps=0
M1016 D_Flip_Flop_5/NAND_0/DS REG_OUT6 gnd Gnd nfet w=8 l=2
+  ad=96 pd=40 as=0 ps=0
M1017 D_Flip_Flop_5/NAND_1/IN_A D_Flip_Flop_3/CLK D_Flip_Flop_5/NAND_0/DS Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1018 D_Flip_Flop_6/QBAR REG_OUT6 vdd vdd pfet w=16 l=2
+  ad=192 pd=56 as=0 ps=0
M1019 vdd D_Flip_Flop_6/NAND_3/IN_B D_Flip_Flop_6/QBAR vdd pfet w=16 l=2
+  ad=0 pd=0 as=0 ps=0
M1020 D_Flip_Flop_6/NAND_3/DS REG_OUT6 gnd Gnd nfet w=8 l=2
+  ad=96 pd=40 as=0 ps=0
M1021 D_Flip_Flop_6/QBAR D_Flip_Flop_6/NAND_3/IN_B D_Flip_Flop_6/NAND_3/DS Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1022 D_Flip_Flop_6/NAND_3/IN_B D_Flip_Flop_6/NAND_2/IN_A vdd vdd pfet w=16 l=2
+  ad=192 pd=56 as=0 ps=0
M1023 vdd D_Flip_Flop_3/CLK D_Flip_Flop_6/NAND_3/IN_B vdd pfet w=16 l=2
+  ad=0 pd=0 as=0 ps=0
M1024 D_Flip_Flop_6/NAND_2/DS D_Flip_Flop_6/NAND_2/IN_A gnd Gnd nfet w=8 l=2
+  ad=96 pd=40 as=0 ps=0
M1025 D_Flip_Flop_6/NAND_3/IN_B D_Flip_Flop_3/CLK D_Flip_Flop_6/NAND_2/DS Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1026 D_Flip_Flop_6/NAND_2/IN_A REG_OUT5 vdd vdd pfet w=16 l=2
+  ad=144 pd=50 as=0 ps=0
M1027 D_Flip_Flop_6/NAND_2/IN_A REG_OUT5 gnd Gnd nfet w=8 l=2
+  ad=72 pd=34 as=0 ps=0
M1028 D_Flip_Flop_6/NAND_1/NAND_AB D_Flip_Flop_6/NAND_1/IN_A vdd vdd pfet w=16 l=2
+  ad=192 pd=56 as=0 ps=0
M1029 vdd D_Flip_Flop_6/QBAR D_Flip_Flop_6/NAND_1/NAND_AB vdd pfet w=16 l=2
+  ad=0 pd=0 as=0 ps=0
M1030 D_Flip_Flop_6/NAND_1/DS D_Flip_Flop_6/NAND_1/IN_A gnd Gnd nfet w=8 l=2
+  ad=96 pd=40 as=0 ps=0
M1031 D_Flip_Flop_6/NAND_1/NAND_AB D_Flip_Flop_6/QBAR D_Flip_Flop_6/NAND_1/DS Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1032 D_Flip_Flop_6/NAND_1/IN_A REG_OUT5 vdd vdd pfet w=16 l=2
+  ad=192 pd=56 as=0 ps=0
M1033 vdd D_Flip_Flop_3/CLK D_Flip_Flop_6/NAND_1/IN_A vdd pfet w=16 l=2
+  ad=0 pd=0 as=0 ps=0
M1034 D_Flip_Flop_6/NAND_0/DS REG_OUT5 gnd Gnd nfet w=8 l=2
+  ad=96 pd=40 as=0 ps=0
M1035 D_Flip_Flop_6/NAND_1/IN_A D_Flip_Flop_3/CLK D_Flip_Flop_6/NAND_0/DS Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1036 D_Flip_Flop_7/QBAR REG_OUT5 vdd vdd pfet w=16 l=2
+  ad=192 pd=56 as=0 ps=0
M1037 vdd D_Flip_Flop_7/NAND_3/IN_B D_Flip_Flop_7/QBAR vdd pfet w=16 l=2
+  ad=0 pd=0 as=0 ps=0
M1038 D_Flip_Flop_7/NAND_3/DS REG_OUT5 gnd Gnd nfet w=8 l=2
+  ad=96 pd=40 as=0 ps=0
M1039 D_Flip_Flop_7/QBAR D_Flip_Flop_7/NAND_3/IN_B D_Flip_Flop_7/NAND_3/DS Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1040 D_Flip_Flop_7/NAND_3/IN_B D_Flip_Flop_7/NAND_2/IN_A vdd vdd pfet w=16 l=2
+  ad=192 pd=56 as=0 ps=0
M1041 vdd D_Flip_Flop_3/CLK D_Flip_Flop_7/NAND_3/IN_B vdd pfet w=16 l=2
+  ad=0 pd=0 as=0 ps=0
M1042 D_Flip_Flop_7/NAND_2/DS D_Flip_Flop_7/NAND_2/IN_A gnd Gnd nfet w=8 l=2
+  ad=96 pd=40 as=0 ps=0
M1043 D_Flip_Flop_7/NAND_3/IN_B D_Flip_Flop_3/CLK D_Flip_Flop_7/NAND_2/DS Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1044 D_Flip_Flop_7/NAND_2/IN_A REG_OUT4 vdd vdd pfet w=16 l=2
+  ad=144 pd=50 as=0 ps=0
M1045 D_Flip_Flop_7/NAND_2/IN_A REG_OUT4 gnd Gnd nfet w=8 l=2
+  ad=72 pd=34 as=0 ps=0
M1046 D_Flip_Flop_7/NAND_1/NAND_AB D_Flip_Flop_7/NAND_1/IN_A vdd vdd pfet w=16 l=2
+  ad=192 pd=56 as=0 ps=0
M1047 vdd D_Flip_Flop_7/QBAR D_Flip_Flop_7/NAND_1/NAND_AB vdd pfet w=16 l=2
+  ad=0 pd=0 as=0 ps=0
M1048 D_Flip_Flop_7/NAND_1/DS D_Flip_Flop_7/NAND_1/IN_A gnd Gnd nfet w=8 l=2
+  ad=96 pd=40 as=0 ps=0
M1049 D_Flip_Flop_7/NAND_1/NAND_AB D_Flip_Flop_7/QBAR D_Flip_Flop_7/NAND_1/DS Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1050 D_Flip_Flop_7/NAND_1/IN_A REG_OUT4 vdd vdd pfet w=16 l=2
+  ad=192 pd=56 as=0 ps=0
M1051 vdd D_Flip_Flop_3/CLK D_Flip_Flop_7/NAND_1/IN_A vdd pfet w=16 l=2
+  ad=0 pd=0 as=0 ps=0
M1052 D_Flip_Flop_7/NAND_0/DS REG_OUT4 gnd Gnd nfet w=8 l=2
+  ad=96 pd=40 as=0 ps=0
M1053 D_Flip_Flop_7/NAND_1/IN_A D_Flip_Flop_3/CLK D_Flip_Flop_7/NAND_0/DS Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1054 D_Flip_Flop_4/QBAR REG_OUT4 vdd vdd pfet w=16 l=2
+  ad=192 pd=56 as=0 ps=0
M1055 vdd D_Flip_Flop_4/NAND_3/IN_B D_Flip_Flop_4/QBAR vdd pfet w=16 l=2
+  ad=0 pd=0 as=0 ps=0
M1056 D_Flip_Flop_4/NAND_3/DS REG_OUT4 gnd Gnd nfet w=8 l=2
+  ad=96 pd=40 as=0 ps=0
M1057 D_Flip_Flop_4/QBAR D_Flip_Flop_4/NAND_3/IN_B D_Flip_Flop_4/NAND_3/DS Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1058 D_Flip_Flop_4/NAND_3/IN_B D_Flip_Flop_4/NAND_2/IN_A vdd vdd pfet w=16 l=2
+  ad=192 pd=56 as=0 ps=0
M1059 vdd D_Flip_Flop_3/CLK D_Flip_Flop_4/NAND_3/IN_B vdd pfet w=16 l=2
+  ad=0 pd=0 as=0 ps=0
M1060 D_Flip_Flop_4/NAND_2/DS D_Flip_Flop_4/NAND_2/IN_A gnd Gnd nfet w=8 l=2
+  ad=96 pd=40 as=0 ps=0
M1061 D_Flip_Flop_4/NAND_3/IN_B D_Flip_Flop_3/CLK D_Flip_Flop_4/NAND_2/DS Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1062 D_Flip_Flop_4/NAND_2/IN_A REG_OUT3 vdd vdd pfet w=16 l=2
+  ad=144 pd=50 as=0 ps=0
M1063 D_Flip_Flop_4/NAND_2/IN_A REG_OUT3 gnd Gnd nfet w=8 l=2
+  ad=72 pd=34 as=0 ps=0
M1064 D_Flip_Flop_4/NAND_1/NAND_AB D_Flip_Flop_4/NAND_1/IN_A vdd vdd pfet w=16 l=2
+  ad=192 pd=56 as=0 ps=0
M1065 vdd D_Flip_Flop_4/QBAR D_Flip_Flop_4/NAND_1/NAND_AB vdd pfet w=16 l=2
+  ad=0 pd=0 as=0 ps=0
M1066 D_Flip_Flop_4/NAND_1/DS D_Flip_Flop_4/NAND_1/IN_A gnd Gnd nfet w=8 l=2
+  ad=96 pd=40 as=0 ps=0
M1067 D_Flip_Flop_4/NAND_1/NAND_AB D_Flip_Flop_4/QBAR D_Flip_Flop_4/NAND_1/DS Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1068 D_Flip_Flop_4/NAND_1/IN_A REG_OUT3 vdd vdd pfet w=16 l=2
+  ad=192 pd=56 as=0 ps=0
M1069 vdd D_Flip_Flop_3/CLK D_Flip_Flop_4/NAND_1/IN_A vdd pfet w=16 l=2
+  ad=0 pd=0 as=0 ps=0
M1070 D_Flip_Flop_4/NAND_0/DS REG_OUT3 gnd Gnd nfet w=8 l=2
+  ad=96 pd=40 as=0 ps=0
M1071 D_Flip_Flop_4/NAND_1/IN_A D_Flip_Flop_3/CLK D_Flip_Flop_4/NAND_0/DS Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1072 D_Flip_Flop_2/QBAR REG_OUT3 vdd vdd pfet w=16 l=2
+  ad=192 pd=56 as=0 ps=0
M1073 vdd D_Flip_Flop_2/NAND_3/IN_B D_Flip_Flop_2/QBAR vdd pfet w=16 l=2
+  ad=0 pd=0 as=0 ps=0
M1074 D_Flip_Flop_2/NAND_3/DS REG_OUT3 gnd Gnd nfet w=8 l=2
+  ad=96 pd=40 as=0 ps=0
M1075 D_Flip_Flop_2/QBAR D_Flip_Flop_2/NAND_3/IN_B D_Flip_Flop_2/NAND_3/DS Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1076 D_Flip_Flop_2/NAND_3/IN_B D_Flip_Flop_2/NAND_2/IN_A vdd vdd pfet w=16 l=2
+  ad=192 pd=56 as=0 ps=0
M1077 vdd D_Flip_Flop_3/CLK D_Flip_Flop_2/NAND_3/IN_B vdd pfet w=16 l=2
+  ad=0 pd=0 as=0 ps=0
M1078 D_Flip_Flop_2/NAND_2/DS D_Flip_Flop_2/NAND_2/IN_A gnd Gnd nfet w=8 l=2
+  ad=96 pd=40 as=0 ps=0
M1079 D_Flip_Flop_2/NAND_3/IN_B D_Flip_Flop_3/CLK D_Flip_Flop_2/NAND_2/DS Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1080 D_Flip_Flop_2/NAND_2/IN_A REG_OUT2 vdd vdd pfet w=16 l=2
+  ad=144 pd=50 as=0 ps=0
M1081 D_Flip_Flop_2/NAND_2/IN_A REG_OUT2 gnd Gnd nfet w=8 l=2
+  ad=72 pd=34 as=0 ps=0
M1082 D_Flip_Flop_2/NAND_1/NAND_AB D_Flip_Flop_2/NAND_1/IN_A vdd vdd pfet w=16 l=2
+  ad=192 pd=56 as=0 ps=0
M1083 vdd D_Flip_Flop_2/QBAR D_Flip_Flop_2/NAND_1/NAND_AB vdd pfet w=16 l=2
+  ad=0 pd=0 as=0 ps=0
M1084 D_Flip_Flop_2/NAND_1/DS D_Flip_Flop_2/NAND_1/IN_A gnd Gnd nfet w=8 l=2
+  ad=96 pd=40 as=0 ps=0
M1085 D_Flip_Flop_2/NAND_1/NAND_AB D_Flip_Flop_2/QBAR D_Flip_Flop_2/NAND_1/DS Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1086 D_Flip_Flop_2/NAND_1/IN_A REG_OUT2 vdd vdd pfet w=16 l=2
+  ad=192 pd=56 as=0 ps=0
M1087 vdd D_Flip_Flop_3/CLK D_Flip_Flop_2/NAND_1/IN_A vdd pfet w=16 l=2
+  ad=0 pd=0 as=0 ps=0
M1088 D_Flip_Flop_2/NAND_0/DS REG_OUT2 gnd Gnd nfet w=8 l=2
+  ad=96 pd=40 as=0 ps=0
M1089 D_Flip_Flop_2/NAND_1/IN_A D_Flip_Flop_3/CLK D_Flip_Flop_2/NAND_0/DS Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1090 D_Flip_Flop_1/QBAR REG_OUT2 vdd vdd pfet w=16 l=2
+  ad=192 pd=56 as=0 ps=0
M1091 vdd D_Flip_Flop_1/NAND_3/IN_B D_Flip_Flop_1/QBAR vdd pfet w=16 l=2
+  ad=0 pd=0 as=0 ps=0
M1092 D_Flip_Flop_1/NAND_3/DS REG_OUT2 gnd Gnd nfet w=8 l=2
+  ad=96 pd=40 as=0 ps=0
M1093 D_Flip_Flop_1/QBAR D_Flip_Flop_1/NAND_3/IN_B D_Flip_Flop_1/NAND_3/DS Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1094 D_Flip_Flop_1/NAND_3/IN_B D_Flip_Flop_1/NAND_2/IN_A vdd vdd pfet w=16 l=2
+  ad=192 pd=56 as=0 ps=0
M1095 vdd D_Flip_Flop_3/CLK D_Flip_Flop_1/NAND_3/IN_B vdd pfet w=16 l=2
+  ad=0 pd=0 as=0 ps=0
M1096 D_Flip_Flop_1/NAND_2/DS D_Flip_Flop_1/NAND_2/IN_A gnd Gnd nfet w=8 l=2
+  ad=96 pd=40 as=0 ps=0
M1097 D_Flip_Flop_1/NAND_3/IN_B D_Flip_Flop_3/CLK D_Flip_Flop_1/NAND_2/DS Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1098 D_Flip_Flop_1/NAND_2/IN_A REG_OUT1 vdd vdd pfet w=16 l=2
+  ad=144 pd=50 as=0 ps=0
M1099 D_Flip_Flop_1/NAND_2/IN_A REG_OUT1 gnd Gnd nfet w=8 l=2
+  ad=72 pd=34 as=0 ps=0
M1100 D_Flip_Flop_1/NAND_1/NAND_AB D_Flip_Flop_1/NAND_1/IN_A vdd vdd pfet w=16 l=2
+  ad=192 pd=56 as=0 ps=0
M1101 vdd D_Flip_Flop_1/QBAR D_Flip_Flop_1/NAND_1/NAND_AB vdd pfet w=16 l=2
+  ad=0 pd=0 as=0 ps=0
M1102 D_Flip_Flop_1/NAND_1/DS D_Flip_Flop_1/NAND_1/IN_A gnd Gnd nfet w=8 l=2
+  ad=96 pd=40 as=0 ps=0
M1103 D_Flip_Flop_1/NAND_1/NAND_AB D_Flip_Flop_1/QBAR D_Flip_Flop_1/NAND_1/DS Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1104 D_Flip_Flop_1/NAND_1/IN_A REG_OUT1 vdd vdd pfet w=16 l=2
+  ad=192 pd=56 as=0 ps=0
M1105 vdd D_Flip_Flop_3/CLK D_Flip_Flop_1/NAND_1/IN_A vdd pfet w=16 l=2
+  ad=0 pd=0 as=0 ps=0
M1106 D_Flip_Flop_1/NAND_0/DS REG_OUT1 gnd Gnd nfet w=8 l=2
+  ad=96 pd=40 as=0 ps=0
M1107 D_Flip_Flop_1/NAND_1/IN_A D_Flip_Flop_3/CLK D_Flip_Flop_1/NAND_0/DS Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1108 D_Flip_Flop_0/QBAR REG_OUT1 vdd vdd pfet w=16 l=2
+  ad=192 pd=56 as=0 ps=0
M1109 vdd D_Flip_Flop_0/NAND_3/IN_B D_Flip_Flop_0/QBAR vdd pfet w=16 l=2
+  ad=0 pd=0 as=0 ps=0
M1110 D_Flip_Flop_0/NAND_3/DS REG_OUT1 gnd Gnd nfet w=8 l=2
+  ad=96 pd=40 as=0 ps=0
M1111 D_Flip_Flop_0/QBAR D_Flip_Flop_0/NAND_3/IN_B D_Flip_Flop_0/NAND_3/DS Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1112 D_Flip_Flop_0/NAND_3/IN_B D_Flip_Flop_0/NAND_2/IN_A vdd vdd pfet w=16 l=2
+  ad=192 pd=56 as=0 ps=0
M1113 vdd D_Flip_Flop_3/CLK D_Flip_Flop_0/NAND_3/IN_B vdd pfet w=16 l=2
+  ad=0 pd=0 as=0 ps=0
M1114 D_Flip_Flop_0/NAND_2/DS D_Flip_Flop_0/NAND_2/IN_A gnd Gnd nfet w=8 l=2
+  ad=96 pd=40 as=0 ps=0
M1115 D_Flip_Flop_0/NAND_3/IN_B D_Flip_Flop_3/CLK D_Flip_Flop_0/NAND_2/DS Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1116 D_Flip_Flop_0/NAND_2/IN_A REG_OUT0 vdd vdd pfet w=16 l=2
+  ad=144 pd=50 as=0 ps=0
M1117 D_Flip_Flop_0/NAND_2/IN_A REG_OUT0 gnd Gnd nfet w=8 l=2
+  ad=72 pd=34 as=0 ps=0
M1118 D_Flip_Flop_0/NAND_1/NAND_AB D_Flip_Flop_0/NAND_1/IN_A vdd vdd pfet w=16 l=2
+  ad=192 pd=56 as=0 ps=0
M1119 vdd D_Flip_Flop_0/QBAR D_Flip_Flop_0/NAND_1/NAND_AB vdd pfet w=16 l=2
+  ad=0 pd=0 as=0 ps=0
M1120 D_Flip_Flop_0/NAND_1/DS D_Flip_Flop_0/NAND_1/IN_A gnd Gnd nfet w=8 l=2
+  ad=96 pd=40 as=0 ps=0
M1121 D_Flip_Flop_0/NAND_1/NAND_AB D_Flip_Flop_0/QBAR D_Flip_Flop_0/NAND_1/DS Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1122 D_Flip_Flop_0/NAND_1/IN_A REG_OUT0 vdd vdd pfet w=16 l=2
+  ad=192 pd=56 as=0 ps=0
M1123 vdd D_Flip_Flop_3/CLK D_Flip_Flop_0/NAND_1/IN_A vdd pfet w=16 l=2
+  ad=0 pd=0 as=0 ps=0
M1124 D_Flip_Flop_0/NAND_0/DS REG_OUT0 gnd Gnd nfet w=8 l=2
+  ad=96 pd=40 as=0 ps=0
M1125 D_Flip_Flop_0/NAND_1/IN_A D_Flip_Flop_3/CLK D_Flip_Flop_0/NAND_0/DS Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1126 D_Flip_Flop_3/QBAR REG_OUT0 vdd vdd pfet w=16 l=2
+  ad=192 pd=56 as=0 ps=0
M1127 vdd D_Flip_Flop_3/NAND_3/IN_B D_Flip_Flop_3/QBAR vdd pfet w=16 l=2
+  ad=0 pd=0 as=0 ps=0
M1128 D_Flip_Flop_3/NAND_3/DS REG_OUT0 gnd Gnd nfet w=8 l=2
+  ad=96 pd=40 as=0 ps=0
M1129 D_Flip_Flop_3/QBAR D_Flip_Flop_3/NAND_3/IN_B D_Flip_Flop_3/NAND_3/DS Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1130 D_Flip_Flop_3/NAND_3/IN_B D_Flip_Flop_3/NAND_2/IN_A vdd vdd pfet w=16 l=2
+  ad=192 pd=56 as=0 ps=0
M1131 vdd D_Flip_Flop_3/CLK D_Flip_Flop_3/NAND_3/IN_B vdd pfet w=16 l=2
+  ad=0 pd=0 as=0 ps=0
M1132 D_Flip_Flop_3/NAND_2/DS D_Flip_Flop_3/NAND_2/IN_A gnd Gnd nfet w=8 l=2
+  ad=96 pd=40 as=0 ps=0
M1133 D_Flip_Flop_3/NAND_3/IN_B D_Flip_Flop_3/CLK D_Flip_Flop_3/NAND_2/DS Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1134 D_Flip_Flop_3/NAND_2/IN_A D_Flip_Flop_3/D vdd vdd pfet w=16 l=2
+  ad=144 pd=50 as=0 ps=0
M1135 D_Flip_Flop_3/NAND_2/IN_A D_Flip_Flop_3/D gnd Gnd nfet w=8 l=2
+  ad=72 pd=34 as=0 ps=0
M1136 D_Flip_Flop_3/NAND_1/NAND_AB D_Flip_Flop_3/NAND_1/IN_A vdd vdd pfet w=16 l=2
+  ad=192 pd=56 as=0 ps=0
M1137 vdd D_Flip_Flop_3/QBAR D_Flip_Flop_3/NAND_1/NAND_AB vdd pfet w=16 l=2
+  ad=0 pd=0 as=0 ps=0
M1138 D_Flip_Flop_3/NAND_1/DS D_Flip_Flop_3/NAND_1/IN_A gnd Gnd nfet w=8 l=2
+  ad=96 pd=40 as=0 ps=0
M1139 D_Flip_Flop_3/NAND_1/NAND_AB D_Flip_Flop_3/QBAR D_Flip_Flop_3/NAND_1/DS Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1140 D_Flip_Flop_3/NAND_1/IN_A D_Flip_Flop_3/D vdd vdd pfet w=16 l=2
+  ad=192 pd=56 as=0 ps=0
M1141 vdd D_Flip_Flop_3/CLK D_Flip_Flop_3/NAND_1/IN_A vdd pfet w=16 l=2
+  ad=0 pd=0 as=0 ps=0
M1142 D_Flip_Flop_3/NAND_0/DS D_Flip_Flop_3/D gnd Gnd nfet w=8 l=2
+  ad=96 pd=40 as=0 ps=0
M1143 D_Flip_Flop_3/NAND_1/IN_A D_Flip_Flop_3/CLK D_Flip_Flop_3/NAND_0/DS Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
C0 vdd D_Flip_Flop_2/QBAR 2.0fF
C1 vdd D_Flip_Flop_4/NAND_1/IN_A 2.0fF
C2 vdd D_Flip_Flop_6/NAND_1/IN_A 2.0fF
C3 vdd D_Flip_Flop_0/QBAR 2.0fF
C4 vdd D_Flip_Flop_3/NAND_3/IN_B 2.0fF
C5 REG_OUT2 vdd 30.4fF
C6 vdd REG_OUT3 30.4fF
C7 vdd D_Flip_Flop_7/NAND_1/IN_A 2.0fF
C8 vdd D_Flip_Flop_3/QBAR 2.0fF
C9 REG_OUT1 vdd 30.4fF
C10 vdd D_Flip_Flop_3/CLK 104.5fF
C11 vdd D_Flip_Flop_2/NAND_1/IN_A 2.0fF
C12 vdd D_Flip_Flop_4/NAND_3/IN_B 2.0fF
C13 D_Flip_Flop_4/QBAR vdd 2.0fF
C14 vdd D_Flip_Flop_5/NAND_1/IN_A 2.0fF
C15 vdd REG_OUT5 30.4fF
C16 REG_OUT7 vdd 2.8fF
C17 vdd D_Flip_Flop_6/QBAR 2.0fF
C18 vdd D_Flip_Flop_5/NAND_3/IN_B 2.0fF
C19 vdd D_Flip_Flop_7/QBAR 2.0fF
C20 vdd D_Flip_Flop_5/QBAR 2.0fF
C21 D_Flip_Flop_3/D vdd 11.3fF
C22 vdd D_Flip_Flop_1/NAND_3/IN_B 2.0fF
C23 vdd D_Flip_Flop_3/NAND_1/IN_A 2.0fF
C24 vdd REG_OUT6 30.4fF
C25 vdd D_Flip_Flop_2/NAND_3/IN_B 2.0fF
C26 vdd REG_OUT4 30.4fF
C27 D_Flip_Flop_1/NAND_1/IN_A vdd 2.0fF
C28 vdd D_Flip_Flop_0/NAND_1/IN_A 2.0fF
C29 vdd REG_OUT0 33.5fF
C30 vdd D_Flip_Flop_0/NAND_3/IN_B 2.0fF
C31 vdd D_Flip_Flop_6/NAND_3/IN_B 2.0fF
C32 vdd D_Flip_Flop_1/QBAR 2.0fF
C33 D_Flip_Flop_7/NAND_3/IN_B vdd 2.0fF
C34 m2_162_18# gnd! 2.7fF **FLOATING
C35 m2_n65_17# gnd! 2.7fF **FLOATING
C36 D_Flip_Flop_3/D gnd! 42.9fF
C37 D_Flip_Flop_3/NAND_1/NAND_AB gnd! 5.3fF
C38 D_Flip_Flop_3/QBAR gnd! 41.9fF
C39 D_Flip_Flop_3/NAND_1/IN_A gnd! 12.8fF
C40 D_Flip_Flop_3/NAND_2/IN_A gnd! 13.1fF
C41 D_Flip_Flop_3/NAND_3/IN_B gnd! 35.2fF
C42 REG_OUT0 gnd! 98.6fF
C43 D_Flip_Flop_0/NAND_1/NAND_AB gnd! 5.3fF
C44 D_Flip_Flop_0/QBAR gnd! 41.9fF
C45 D_Flip_Flop_0/NAND_1/IN_A gnd! 12.8fF
C46 D_Flip_Flop_0/NAND_2/IN_A gnd! 13.1fF
C47 D_Flip_Flop_0/NAND_3/IN_B gnd! 35.2fF
C48 REG_OUT1 gnd! 98.8fF
C49 D_Flip_Flop_1/NAND_1/NAND_AB gnd! 5.3fF
C50 D_Flip_Flop_1/QBAR gnd! 41.9fF
C51 D_Flip_Flop_1/NAND_1/IN_A gnd! 12.8fF
C52 D_Flip_Flop_1/NAND_2/IN_A gnd! 13.1fF
C53 D_Flip_Flop_1/NAND_3/IN_B gnd! 35.2fF
C54 REG_OUT2 gnd! 98.7fF
C55 D_Flip_Flop_2/NAND_1/NAND_AB gnd! 5.3fF
C56 D_Flip_Flop_2/QBAR gnd! 41.9fF
C57 D_Flip_Flop_2/NAND_1/IN_A gnd! 12.8fF
C58 D_Flip_Flop_2/NAND_2/IN_A gnd! 13.1fF
C59 D_Flip_Flop_2/NAND_3/IN_B gnd! 35.2fF
C60 REG_OUT3 gnd! 96.5fF
C61 D_Flip_Flop_4/NAND_1/NAND_AB gnd! 5.3fF
C62 D_Flip_Flop_4/QBAR gnd! 41.9fF
C63 D_Flip_Flop_4/NAND_1/IN_A gnd! 12.8fF
C64 D_Flip_Flop_4/NAND_2/IN_A gnd! 13.1fF
C65 D_Flip_Flop_4/NAND_3/IN_B gnd! 35.2fF
C66 REG_OUT4 gnd! 99.1fF
C67 D_Flip_Flop_7/NAND_1/NAND_AB gnd! 5.3fF
C68 D_Flip_Flop_7/QBAR gnd! 41.9fF
C69 D_Flip_Flop_7/NAND_1/IN_A gnd! 12.8fF
C70 D_Flip_Flop_7/NAND_2/IN_A gnd! 13.1fF
C71 D_Flip_Flop_7/NAND_3/IN_B gnd! 35.2fF
C72 REG_OUT5 gnd! 98.8fF
C73 D_Flip_Flop_6/NAND_1/NAND_AB gnd! 5.3fF
C74 D_Flip_Flop_6/QBAR gnd! 41.9fF
C75 D_Flip_Flop_6/NAND_1/IN_A gnd! 12.8fF
C76 D_Flip_Flop_6/NAND_2/IN_A gnd! 13.1fF
C77 D_Flip_Flop_6/NAND_3/IN_B gnd! 35.2fF
C78 D_Flip_Flop_3/CLK gnd! 1133.0fF
C79 REG_OUT6 gnd! 97.8fF
C80 D_Flip_Flop_5/NAND_1/NAND_AB gnd! 5.3fF
C81 D_Flip_Flop_5/QBAR gnd! 41.9fF
C82 D_Flip_Flop_5/NAND_1/IN_A gnd! 12.8fF
C83 vdd gnd! 4215.9fF
C84 D_Flip_Flop_5/NAND_2/IN_A gnd! 13.1fF
C85 D_Flip_Flop_5/NAND_3/IN_B gnd! 35.2fF
C86 REG_OUT7 gnd! 60.2fF
