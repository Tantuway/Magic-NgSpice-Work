* SPICE3 file created from 8BITadder.ext - technology: scmos

.option scale=1u

M1000 FULL_ADDER_7/COUT FULL_ADDER_7/NAND_2/IN_A vdd vdd pfet w=16 l=2
+  ad=192 pd=56 as=9472 ps=4768
M1001 vdd FULL_ADDER_7/NAND_2/IN_B FULL_ADDER_7/COUT vdd pfet w=16 l=2
+  ad=0 pd=0 as=0 ps=0
M1002 FULL_ADDER_7/NAND_2/DS FULL_ADDER_7/NAND_2/IN_A gnd Gnd nfet w=8 l=2
+  ad=96 pd=40 as=3520 ps=2288
M1003 FULL_ADDER_7/COUT FULL_ADDER_7/NAND_2/IN_B FULL_ADDER_7/NAND_2/DS Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1004 FULL_ADDER_7/NAND_2/IN_B FULL_ADDER_7/B vdd vdd pfet w=16 l=2
+  ad=192 pd=56 as=0 ps=0
M1005 vdd gnd FULL_ADDER_7/NAND_2/IN_B vdd pfet w=16 l=2
+  ad=0 pd=0 as=0 ps=0
M1006 FULL_ADDER_7/NAND_1/DS FULL_ADDER_7/B gnd Gnd nfet w=8 l=2
+  ad=96 pd=40 as=0 ps=0
M1007 FULL_ADDER_7/NAND_2/IN_B gnd FULL_ADDER_7/NAND_1/DS Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1008 FULL_ADDER_7/NAND_2/IN_A FULL_ADDER_7/CIN vdd vdd pfet w=16 l=2
+  ad=192 pd=56 as=0 ps=0
M1009 vdd FULL_ADDER_7/XOR_1/A FULL_ADDER_7/NAND_2/IN_A vdd pfet w=16 l=2
+  ad=0 pd=0 as=0 ps=0
M1010 FULL_ADDER_7/NAND_0/DS FULL_ADDER_7/CIN gnd Gnd nfet w=8 l=2
+  ad=96 pd=40 as=0 ps=0
M1011 FULL_ADDER_7/NAND_2/IN_A FULL_ADDER_7/XOR_1/A FULL_ADDER_7/NAND_0/DS Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1012 FULL_ADDER_7/XOR_1/a_n3_n2# FULL_ADDER_7/XOR_1/A vdd FULL_ADDER_7/XOR_1/w_n16_50# pfet w=16 l=2
+  ad=96 pd=44 as=0 ps=0
M1013 FULL_ADDER_7/XOR_1/a_18_52# FULL_ADDER_7/XOR_1/a_n3_n2# vdd FULL_ADDER_7/XOR_1/w_n16_50# pfet w=16 l=2
+  ad=80 pd=42 as=0 ps=0
M1014 FULL_ADDER_7/SUM FULL_ADDER_7/CIN FULL_ADDER_7/XOR_1/a_18_52# FULL_ADDER_7/XOR_1/w_n16_50# pfet w=16 l=2
+  ad=224 pd=92 as=0 ps=0
M1015 FULL_ADDER_7/XOR_1/a_47_52# FULL_ADDER_7/XOR_1/a_21_19# FULL_ADDER_7/SUM FULL_ADDER_7/XOR_1/w_n16_50# pfet w=16 l=2
+  ad=80 pd=42 as=0 ps=0
M1016 vdd FULL_ADDER_7/XOR_1/a_52_45# FULL_ADDER_7/XOR_1/a_47_52# FULL_ADDER_7/XOR_1/w_n16_50# pfet w=16 l=2
+  ad=0 pd=0 as=0 ps=0
M1017 vdd FULL_ADDER_7/CIN FULL_ADDER_7/XOR_1/a_52_45# FULL_ADDER_7/XOR_1/w_n16_50# pfet w=16 l=2
+  ad=0 pd=0 as=96 ps=44
M1018 FULL_ADDER_7/XOR_1/a_n3_n2# FULL_ADDER_7/XOR_1/A gnd Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1019 FULL_ADDER_7/XOR_1/a_18_n2# FULL_ADDER_7/CIN gnd Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1020 FULL_ADDER_7/SUM FULL_ADDER_7/XOR_1/a_21_19# FULL_ADDER_7/XOR_1/a_18_n2# Gnd nfet w=8 l=2
+  ad=120 pd=62 as=0 ps=0
M1021 FULL_ADDER_7/XOR_1/a_48_n2# FULL_ADDER_7/XOR_1/a_n3_n2# FULL_ADDER_7/SUM Gnd nfet w=8 l=2
+  ad=48 pd=28 as=0 ps=0
M1022 gnd FULL_ADDER_7/XOR_1/a_52_45# FULL_ADDER_7/XOR_1/a_48_n2# Gnd nfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1023 gnd FULL_ADDER_7/CIN FULL_ADDER_7/XOR_1/a_52_45# Gnd nfet w=8 l=2
+  ad=0 pd=0 as=40 ps=26
M1024 FULL_ADDER_7/XOR_0/a_n3_n2# FULL_ADDER_7/XOR_0/A vdd FULL_ADDER_7/XOR_0/w_n16_50# pfet w=16 l=2
+  ad=96 pd=44 as=0 ps=0
M1025 FULL_ADDER_7/XOR_0/a_18_52# FULL_ADDER_7/XOR_0/a_n3_n2# vdd FULL_ADDER_7/XOR_0/w_n16_50# pfet w=16 l=2
+  ad=80 pd=42 as=0 ps=0
M1026 FULL_ADDER_7/XOR_1/A FULL_ADDER_7/B FULL_ADDER_7/XOR_0/a_18_52# FULL_ADDER_7/XOR_0/w_n16_50# pfet w=16 l=2
+  ad=224 pd=92 as=0 ps=0
M1027 FULL_ADDER_7/XOR_0/a_47_52# FULL_ADDER_7/XOR_0/a_21_19# FULL_ADDER_7/XOR_1/A FULL_ADDER_7/XOR_0/w_n16_50# pfet w=16 l=2
+  ad=80 pd=42 as=0 ps=0
M1028 vdd FULL_ADDER_7/XOR_0/a_52_45# FULL_ADDER_7/XOR_0/a_47_52# FULL_ADDER_7/XOR_0/w_n16_50# pfet w=16 l=2
+  ad=0 pd=0 as=0 ps=0
M1029 vdd FULL_ADDER_7/B FULL_ADDER_7/XOR_0/a_52_45# FULL_ADDER_7/XOR_0/w_n16_50# pfet w=16 l=2
+  ad=0 pd=0 as=96 ps=44
M1030 FULL_ADDER_7/XOR_0/a_n3_n2# FULL_ADDER_7/XOR_0/A gnd Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1031 FULL_ADDER_7/XOR_0/a_18_n2# FULL_ADDER_7/B gnd Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1032 FULL_ADDER_7/XOR_1/A FULL_ADDER_7/XOR_0/a_21_19# FULL_ADDER_7/XOR_0/a_18_n2# Gnd nfet w=8 l=2
+  ad=120 pd=62 as=0 ps=0
M1033 FULL_ADDER_7/XOR_0/a_48_n2# FULL_ADDER_7/XOR_0/a_n3_n2# FULL_ADDER_7/XOR_1/A Gnd nfet w=8 l=2
+  ad=48 pd=28 as=0 ps=0
M1034 gnd FULL_ADDER_7/XOR_0/a_52_45# FULL_ADDER_7/XOR_0/a_48_n2# Gnd nfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1035 gnd FULL_ADDER_7/B FULL_ADDER_7/XOR_0/a_52_45# Gnd nfet w=8 l=2
+  ad=0 pd=0 as=40 ps=26
M1036 FULL_ADDER_6/COUT FULL_ADDER_6/NAND_2/IN_A vdd vdd pfet w=16 l=2
+  ad=192 pd=56 as=0 ps=0
M1037 vdd FULL_ADDER_6/NAND_2/IN_B FULL_ADDER_6/COUT vdd pfet w=16 l=2
+  ad=0 pd=0 as=0 ps=0
M1038 FULL_ADDER_6/NAND_2/DS FULL_ADDER_6/NAND_2/IN_A gnd Gnd nfet w=8 l=2
+  ad=96 pd=40 as=0 ps=0
M1039 FULL_ADDER_6/COUT FULL_ADDER_6/NAND_2/IN_B FULL_ADDER_6/NAND_2/DS Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1040 FULL_ADDER_6/NAND_2/IN_B FULL_ADDER_6/B vdd vdd pfet w=16 l=2
+  ad=192 pd=56 as=0 ps=0
M1041 vdd gnd FULL_ADDER_6/NAND_2/IN_B vdd pfet w=16 l=2
+  ad=0 pd=0 as=0 ps=0
M1042 FULL_ADDER_6/NAND_1/DS FULL_ADDER_6/B gnd Gnd nfet w=8 l=2
+  ad=96 pd=40 as=0 ps=0
M1043 FULL_ADDER_6/NAND_2/IN_B gnd FULL_ADDER_6/NAND_1/DS Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1044 FULL_ADDER_6/NAND_2/IN_A FULL_ADDER_6/CIN vdd vdd pfet w=16 l=2
+  ad=192 pd=56 as=0 ps=0
M1045 vdd FULL_ADDER_6/XOR_1/A FULL_ADDER_6/NAND_2/IN_A vdd pfet w=16 l=2
+  ad=0 pd=0 as=0 ps=0
M1046 FULL_ADDER_6/NAND_0/DS FULL_ADDER_6/CIN gnd Gnd nfet w=8 l=2
+  ad=96 pd=40 as=0 ps=0
M1047 FULL_ADDER_6/NAND_2/IN_A FULL_ADDER_6/XOR_1/A FULL_ADDER_6/NAND_0/DS Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1048 FULL_ADDER_6/XOR_1/a_n3_n2# FULL_ADDER_6/XOR_1/A vdd FULL_ADDER_6/XOR_1/w_n16_50# pfet w=16 l=2
+  ad=96 pd=44 as=0 ps=0
M1049 FULL_ADDER_6/XOR_1/a_18_52# FULL_ADDER_6/XOR_1/a_n3_n2# vdd FULL_ADDER_6/XOR_1/w_n16_50# pfet w=16 l=2
+  ad=80 pd=42 as=0 ps=0
M1050 FULL_ADDER_6/SUM FULL_ADDER_6/CIN FULL_ADDER_6/XOR_1/a_18_52# FULL_ADDER_6/XOR_1/w_n16_50# pfet w=16 l=2
+  ad=224 pd=92 as=0 ps=0
M1051 FULL_ADDER_6/XOR_1/a_47_52# FULL_ADDER_6/XOR_1/a_21_19# FULL_ADDER_6/SUM FULL_ADDER_6/XOR_1/w_n16_50# pfet w=16 l=2
+  ad=80 pd=42 as=0 ps=0
M1052 vdd FULL_ADDER_6/XOR_1/a_52_45# FULL_ADDER_6/XOR_1/a_47_52# FULL_ADDER_6/XOR_1/w_n16_50# pfet w=16 l=2
+  ad=0 pd=0 as=0 ps=0
M1053 vdd FULL_ADDER_6/CIN FULL_ADDER_6/XOR_1/a_52_45# FULL_ADDER_6/XOR_1/w_n16_50# pfet w=16 l=2
+  ad=0 pd=0 as=96 ps=44
M1054 FULL_ADDER_6/XOR_1/a_n3_n2# FULL_ADDER_6/XOR_1/A gnd Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1055 FULL_ADDER_6/XOR_1/a_18_n2# FULL_ADDER_6/CIN gnd Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1056 FULL_ADDER_6/SUM FULL_ADDER_6/XOR_1/a_21_19# FULL_ADDER_6/XOR_1/a_18_n2# Gnd nfet w=8 l=2
+  ad=120 pd=62 as=0 ps=0
M1057 FULL_ADDER_6/XOR_1/a_48_n2# FULL_ADDER_6/XOR_1/a_n3_n2# FULL_ADDER_6/SUM Gnd nfet w=8 l=2
+  ad=48 pd=28 as=0 ps=0
M1058 gnd FULL_ADDER_6/XOR_1/a_52_45# FULL_ADDER_6/XOR_1/a_48_n2# Gnd nfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1059 gnd FULL_ADDER_6/CIN FULL_ADDER_6/XOR_1/a_52_45# Gnd nfet w=8 l=2
+  ad=0 pd=0 as=40 ps=26
M1060 FULL_ADDER_6/XOR_0/a_n3_n2# FULL_ADDER_6/XOR_0/A vdd FULL_ADDER_6/XOR_0/w_n16_50# pfet w=16 l=2
+  ad=96 pd=44 as=0 ps=0
M1061 FULL_ADDER_6/XOR_0/a_18_52# FULL_ADDER_6/XOR_0/a_n3_n2# vdd FULL_ADDER_6/XOR_0/w_n16_50# pfet w=16 l=2
+  ad=80 pd=42 as=0 ps=0
M1062 FULL_ADDER_6/XOR_1/A FULL_ADDER_6/B FULL_ADDER_6/XOR_0/a_18_52# FULL_ADDER_6/XOR_0/w_n16_50# pfet w=16 l=2
+  ad=224 pd=92 as=0 ps=0
M1063 FULL_ADDER_6/XOR_0/a_47_52# FULL_ADDER_6/XOR_0/a_21_19# FULL_ADDER_6/XOR_1/A FULL_ADDER_6/XOR_0/w_n16_50# pfet w=16 l=2
+  ad=80 pd=42 as=0 ps=0
M1064 vdd FULL_ADDER_6/XOR_0/a_52_45# FULL_ADDER_6/XOR_0/a_47_52# FULL_ADDER_6/XOR_0/w_n16_50# pfet w=16 l=2
+  ad=0 pd=0 as=0 ps=0
M1065 vdd FULL_ADDER_6/B FULL_ADDER_6/XOR_0/a_52_45# FULL_ADDER_6/XOR_0/w_n16_50# pfet w=16 l=2
+  ad=0 pd=0 as=96 ps=44
M1066 FULL_ADDER_6/XOR_0/a_n3_n2# FULL_ADDER_6/XOR_0/A gnd Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1067 FULL_ADDER_6/XOR_0/a_18_n2# FULL_ADDER_6/B gnd Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1068 FULL_ADDER_6/XOR_1/A FULL_ADDER_6/XOR_0/a_21_19# FULL_ADDER_6/XOR_0/a_18_n2# Gnd nfet w=8 l=2
+  ad=120 pd=62 as=0 ps=0
M1069 FULL_ADDER_6/XOR_0/a_48_n2# FULL_ADDER_6/XOR_0/a_n3_n2# FULL_ADDER_6/XOR_1/A Gnd nfet w=8 l=2
+  ad=48 pd=28 as=0 ps=0
M1070 gnd FULL_ADDER_6/XOR_0/a_52_45# FULL_ADDER_6/XOR_0/a_48_n2# Gnd nfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1071 gnd FULL_ADDER_6/B FULL_ADDER_6/XOR_0/a_52_45# Gnd nfet w=8 l=2
+  ad=0 pd=0 as=40 ps=26
M1072 FULL_ADDER_5/COUT FULL_ADDER_5/NAND_2/IN_A vdd vdd pfet w=16 l=2
+  ad=192 pd=56 as=0 ps=0
M1073 vdd FULL_ADDER_5/NAND_2/IN_B FULL_ADDER_5/COUT vdd pfet w=16 l=2
+  ad=0 pd=0 as=0 ps=0
M1074 FULL_ADDER_5/NAND_2/DS FULL_ADDER_5/NAND_2/IN_A gnd Gnd nfet w=8 l=2
+  ad=96 pd=40 as=0 ps=0
M1075 FULL_ADDER_5/COUT FULL_ADDER_5/NAND_2/IN_B FULL_ADDER_5/NAND_2/DS Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1076 FULL_ADDER_5/NAND_2/IN_B FULL_ADDER_5/B vdd vdd pfet w=16 l=2
+  ad=192 pd=56 as=0 ps=0
M1077 vdd gnd FULL_ADDER_5/NAND_2/IN_B vdd pfet w=16 l=2
+  ad=0 pd=0 as=0 ps=0
M1078 FULL_ADDER_5/NAND_1/DS FULL_ADDER_5/B gnd Gnd nfet w=8 l=2
+  ad=96 pd=40 as=0 ps=0
M1079 FULL_ADDER_5/NAND_2/IN_B gnd FULL_ADDER_5/NAND_1/DS Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1080 FULL_ADDER_5/NAND_2/IN_A FULL_ADDER_5/CIN vdd vdd pfet w=16 l=2
+  ad=192 pd=56 as=0 ps=0
M1081 vdd FULL_ADDER_5/XOR_1/A FULL_ADDER_5/NAND_2/IN_A vdd pfet w=16 l=2
+  ad=0 pd=0 as=0 ps=0
M1082 FULL_ADDER_5/NAND_0/DS FULL_ADDER_5/CIN gnd Gnd nfet w=8 l=2
+  ad=96 pd=40 as=0 ps=0
M1083 FULL_ADDER_5/NAND_2/IN_A FULL_ADDER_5/XOR_1/A FULL_ADDER_5/NAND_0/DS Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1084 FULL_ADDER_5/XOR_1/a_n3_n2# FULL_ADDER_5/XOR_1/A vdd FULL_ADDER_5/XOR_1/w_n16_50# pfet w=16 l=2
+  ad=96 pd=44 as=0 ps=0
M1085 FULL_ADDER_5/XOR_1/a_18_52# FULL_ADDER_5/XOR_1/a_n3_n2# vdd FULL_ADDER_5/XOR_1/w_n16_50# pfet w=16 l=2
+  ad=80 pd=42 as=0 ps=0
M1086 FULL_ADDER_5/SUM FULL_ADDER_5/CIN FULL_ADDER_5/XOR_1/a_18_52# FULL_ADDER_5/XOR_1/w_n16_50# pfet w=16 l=2
+  ad=224 pd=92 as=0 ps=0
M1087 FULL_ADDER_5/XOR_1/a_47_52# FULL_ADDER_5/XOR_1/a_21_19# FULL_ADDER_5/SUM FULL_ADDER_5/XOR_1/w_n16_50# pfet w=16 l=2
+  ad=80 pd=42 as=0 ps=0
M1088 vdd FULL_ADDER_5/XOR_1/a_52_45# FULL_ADDER_5/XOR_1/a_47_52# FULL_ADDER_5/XOR_1/w_n16_50# pfet w=16 l=2
+  ad=0 pd=0 as=0 ps=0
M1089 vdd FULL_ADDER_5/CIN FULL_ADDER_5/XOR_1/a_52_45# FULL_ADDER_5/XOR_1/w_n16_50# pfet w=16 l=2
+  ad=0 pd=0 as=96 ps=44
M1090 FULL_ADDER_5/XOR_1/a_n3_n2# FULL_ADDER_5/XOR_1/A gnd Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1091 FULL_ADDER_5/XOR_1/a_18_n2# FULL_ADDER_5/CIN gnd Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1092 FULL_ADDER_5/SUM FULL_ADDER_5/XOR_1/a_21_19# FULL_ADDER_5/XOR_1/a_18_n2# Gnd nfet w=8 l=2
+  ad=120 pd=62 as=0 ps=0
M1093 FULL_ADDER_5/XOR_1/a_48_n2# FULL_ADDER_5/XOR_1/a_n3_n2# FULL_ADDER_5/SUM Gnd nfet w=8 l=2
+  ad=48 pd=28 as=0 ps=0
M1094 gnd FULL_ADDER_5/XOR_1/a_52_45# FULL_ADDER_5/XOR_1/a_48_n2# Gnd nfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1095 gnd FULL_ADDER_5/CIN FULL_ADDER_5/XOR_1/a_52_45# Gnd nfet w=8 l=2
+  ad=0 pd=0 as=40 ps=26
M1096 FULL_ADDER_5/XOR_0/a_n3_n2# FULL_ADDER_5/XOR_0/A vdd FULL_ADDER_5/XOR_0/w_n16_50# pfet w=16 l=2
+  ad=96 pd=44 as=0 ps=0
M1097 FULL_ADDER_5/XOR_0/a_18_52# FULL_ADDER_5/XOR_0/a_n3_n2# vdd FULL_ADDER_5/XOR_0/w_n16_50# pfet w=16 l=2
+  ad=80 pd=42 as=0 ps=0
M1098 FULL_ADDER_5/XOR_1/A FULL_ADDER_5/B FULL_ADDER_5/XOR_0/a_18_52# FULL_ADDER_5/XOR_0/w_n16_50# pfet w=16 l=2
+  ad=224 pd=92 as=0 ps=0
M1099 FULL_ADDER_5/XOR_0/a_47_52# FULL_ADDER_5/XOR_0/a_21_19# FULL_ADDER_5/XOR_1/A FULL_ADDER_5/XOR_0/w_n16_50# pfet w=16 l=2
+  ad=80 pd=42 as=0 ps=0
M1100 vdd FULL_ADDER_5/XOR_0/a_52_45# FULL_ADDER_5/XOR_0/a_47_52# FULL_ADDER_5/XOR_0/w_n16_50# pfet w=16 l=2
+  ad=0 pd=0 as=0 ps=0
M1101 vdd FULL_ADDER_5/B FULL_ADDER_5/XOR_0/a_52_45# FULL_ADDER_5/XOR_0/w_n16_50# pfet w=16 l=2
+  ad=0 pd=0 as=96 ps=44
M1102 FULL_ADDER_5/XOR_0/a_n3_n2# FULL_ADDER_5/XOR_0/A gnd Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1103 FULL_ADDER_5/XOR_0/a_18_n2# FULL_ADDER_5/B gnd Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1104 FULL_ADDER_5/XOR_1/A FULL_ADDER_5/XOR_0/a_21_19# FULL_ADDER_5/XOR_0/a_18_n2# Gnd nfet w=8 l=2
+  ad=120 pd=62 as=0 ps=0
M1105 FULL_ADDER_5/XOR_0/a_48_n2# FULL_ADDER_5/XOR_0/a_n3_n2# FULL_ADDER_5/XOR_1/A Gnd nfet w=8 l=2
+  ad=48 pd=28 as=0 ps=0
M1106 gnd FULL_ADDER_5/XOR_0/a_52_45# FULL_ADDER_5/XOR_0/a_48_n2# Gnd nfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1107 gnd FULL_ADDER_5/B FULL_ADDER_5/XOR_0/a_52_45# Gnd nfet w=8 l=2
+  ad=0 pd=0 as=40 ps=26
M1108 FULL_ADDER_4/COUT FULL_ADDER_4/NAND_2/IN_A vdd vdd pfet w=16 l=2
+  ad=192 pd=56 as=0 ps=0
M1109 vdd FULL_ADDER_4/NAND_2/IN_B FULL_ADDER_4/COUT vdd pfet w=16 l=2
+  ad=0 pd=0 as=0 ps=0
M1110 FULL_ADDER_4/NAND_2/DS FULL_ADDER_4/NAND_2/IN_A gnd Gnd nfet w=8 l=2
+  ad=96 pd=40 as=0 ps=0
M1111 FULL_ADDER_4/COUT FULL_ADDER_4/NAND_2/IN_B FULL_ADDER_4/NAND_2/DS Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1112 FULL_ADDER_4/NAND_2/IN_B FULL_ADDER_4/B vdd vdd pfet w=16 l=2
+  ad=192 pd=56 as=0 ps=0
M1113 vdd gnd FULL_ADDER_4/NAND_2/IN_B vdd pfet w=16 l=2
+  ad=0 pd=0 as=0 ps=0
M1114 FULL_ADDER_4/NAND_1/DS FULL_ADDER_4/B gnd Gnd nfet w=8 l=2
+  ad=96 pd=40 as=0 ps=0
M1115 FULL_ADDER_4/NAND_2/IN_B gnd FULL_ADDER_4/NAND_1/DS Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1116 FULL_ADDER_4/NAND_2/IN_A FULL_ADDER_4/CIN vdd vdd pfet w=16 l=2
+  ad=192 pd=56 as=0 ps=0
M1117 vdd FULL_ADDER_4/XOR_1/A FULL_ADDER_4/NAND_2/IN_A vdd pfet w=16 l=2
+  ad=0 pd=0 as=0 ps=0
M1118 FULL_ADDER_4/NAND_0/DS FULL_ADDER_4/CIN gnd Gnd nfet w=8 l=2
+  ad=96 pd=40 as=0 ps=0
M1119 FULL_ADDER_4/NAND_2/IN_A FULL_ADDER_4/XOR_1/A FULL_ADDER_4/NAND_0/DS Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1120 FULL_ADDER_4/XOR_1/a_n3_n2# FULL_ADDER_4/XOR_1/A vdd FULL_ADDER_4/XOR_1/w_n16_50# pfet w=16 l=2
+  ad=96 pd=44 as=0 ps=0
M1121 FULL_ADDER_4/XOR_1/a_18_52# FULL_ADDER_4/XOR_1/a_n3_n2# vdd FULL_ADDER_4/XOR_1/w_n16_50# pfet w=16 l=2
+  ad=80 pd=42 as=0 ps=0
M1122 FULL_ADDER_4/SUM FULL_ADDER_4/CIN FULL_ADDER_4/XOR_1/a_18_52# FULL_ADDER_4/XOR_1/w_n16_50# pfet w=16 l=2
+  ad=224 pd=92 as=0 ps=0
M1123 FULL_ADDER_4/XOR_1/a_47_52# FULL_ADDER_4/XOR_1/a_21_19# FULL_ADDER_4/SUM FULL_ADDER_4/XOR_1/w_n16_50# pfet w=16 l=2
+  ad=80 pd=42 as=0 ps=0
M1124 vdd FULL_ADDER_4/XOR_1/a_52_45# FULL_ADDER_4/XOR_1/a_47_52# FULL_ADDER_4/XOR_1/w_n16_50# pfet w=16 l=2
+  ad=0 pd=0 as=0 ps=0
M1125 vdd FULL_ADDER_4/CIN FULL_ADDER_4/XOR_1/a_52_45# FULL_ADDER_4/XOR_1/w_n16_50# pfet w=16 l=2
+  ad=0 pd=0 as=96 ps=44
M1126 FULL_ADDER_4/XOR_1/a_n3_n2# FULL_ADDER_4/XOR_1/A gnd Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1127 FULL_ADDER_4/XOR_1/a_18_n2# FULL_ADDER_4/CIN gnd Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1128 FULL_ADDER_4/SUM FULL_ADDER_4/XOR_1/a_21_19# FULL_ADDER_4/XOR_1/a_18_n2# Gnd nfet w=8 l=2
+  ad=120 pd=62 as=0 ps=0
M1129 FULL_ADDER_4/XOR_1/a_48_n2# FULL_ADDER_4/XOR_1/a_n3_n2# FULL_ADDER_4/SUM Gnd nfet w=8 l=2
+  ad=48 pd=28 as=0 ps=0
M1130 gnd FULL_ADDER_4/XOR_1/a_52_45# FULL_ADDER_4/XOR_1/a_48_n2# Gnd nfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1131 gnd FULL_ADDER_4/CIN FULL_ADDER_4/XOR_1/a_52_45# Gnd nfet w=8 l=2
+  ad=0 pd=0 as=40 ps=26
M1132 FULL_ADDER_4/XOR_0/a_n3_n2# FULL_ADDER_4/XOR_0/A vdd FULL_ADDER_4/XOR_0/w_n16_50# pfet w=16 l=2
+  ad=96 pd=44 as=0 ps=0
M1133 FULL_ADDER_4/XOR_0/a_18_52# FULL_ADDER_4/XOR_0/a_n3_n2# vdd FULL_ADDER_4/XOR_0/w_n16_50# pfet w=16 l=2
+  ad=80 pd=42 as=0 ps=0
M1134 FULL_ADDER_4/XOR_1/A FULL_ADDER_4/B FULL_ADDER_4/XOR_0/a_18_52# FULL_ADDER_4/XOR_0/w_n16_50# pfet w=16 l=2
+  ad=224 pd=92 as=0 ps=0
M1135 FULL_ADDER_4/XOR_0/a_47_52# FULL_ADDER_4/XOR_0/a_21_19# FULL_ADDER_4/XOR_1/A FULL_ADDER_4/XOR_0/w_n16_50# pfet w=16 l=2
+  ad=80 pd=42 as=0 ps=0
M1136 vdd FULL_ADDER_4/XOR_0/a_52_45# FULL_ADDER_4/XOR_0/a_47_52# FULL_ADDER_4/XOR_0/w_n16_50# pfet w=16 l=2
+  ad=0 pd=0 as=0 ps=0
M1137 vdd FULL_ADDER_4/B FULL_ADDER_4/XOR_0/a_52_45# FULL_ADDER_4/XOR_0/w_n16_50# pfet w=16 l=2
+  ad=0 pd=0 as=96 ps=44
M1138 FULL_ADDER_4/XOR_0/a_n3_n2# FULL_ADDER_4/XOR_0/A gnd Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1139 FULL_ADDER_4/XOR_0/a_18_n2# FULL_ADDER_4/B gnd Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1140 FULL_ADDER_4/XOR_1/A FULL_ADDER_4/XOR_0/a_21_19# FULL_ADDER_4/XOR_0/a_18_n2# Gnd nfet w=8 l=2
+  ad=120 pd=62 as=0 ps=0
M1141 FULL_ADDER_4/XOR_0/a_48_n2# FULL_ADDER_4/XOR_0/a_n3_n2# FULL_ADDER_4/XOR_1/A Gnd nfet w=8 l=2
+  ad=48 pd=28 as=0 ps=0
M1142 gnd FULL_ADDER_4/XOR_0/a_52_45# FULL_ADDER_4/XOR_0/a_48_n2# Gnd nfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1143 gnd FULL_ADDER_4/B FULL_ADDER_4/XOR_0/a_52_45# Gnd nfet w=8 l=2
+  ad=0 pd=0 as=40 ps=26
M1144 FULL_ADDER_3/COUT FULL_ADDER_3/NAND_2/IN_A vdd vdd pfet w=16 l=2
+  ad=192 pd=56 as=0 ps=0
M1145 vdd FULL_ADDER_3/NAND_2/IN_B FULL_ADDER_3/COUT vdd pfet w=16 l=2
+  ad=0 pd=0 as=0 ps=0
M1146 FULL_ADDER_3/NAND_2/DS FULL_ADDER_3/NAND_2/IN_A gnd Gnd nfet w=8 l=2
+  ad=96 pd=40 as=0 ps=0
M1147 FULL_ADDER_3/COUT FULL_ADDER_3/NAND_2/IN_B FULL_ADDER_3/NAND_2/DS Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1148 FULL_ADDER_3/NAND_2/IN_B FULL_ADDER_3/B vdd vdd pfet w=16 l=2
+  ad=192 pd=56 as=0 ps=0
M1149 vdd gnd FULL_ADDER_3/NAND_2/IN_B vdd pfet w=16 l=2
+  ad=0 pd=0 as=0 ps=0
M1150 FULL_ADDER_3/NAND_1/DS FULL_ADDER_3/B gnd Gnd nfet w=8 l=2
+  ad=96 pd=40 as=0 ps=0
M1151 FULL_ADDER_3/NAND_2/IN_B gnd FULL_ADDER_3/NAND_1/DS Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1152 FULL_ADDER_3/NAND_2/IN_A FULL_ADDER_3/CIN vdd vdd pfet w=16 l=2
+  ad=192 pd=56 as=0 ps=0
M1153 vdd FULL_ADDER_3/XOR_1/A FULL_ADDER_3/NAND_2/IN_A vdd pfet w=16 l=2
+  ad=0 pd=0 as=0 ps=0
M1154 FULL_ADDER_3/NAND_0/DS FULL_ADDER_3/CIN gnd Gnd nfet w=8 l=2
+  ad=96 pd=40 as=0 ps=0
M1155 FULL_ADDER_3/NAND_2/IN_A FULL_ADDER_3/XOR_1/A FULL_ADDER_3/NAND_0/DS Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1156 FULL_ADDER_3/XOR_1/a_n3_n2# FULL_ADDER_3/XOR_1/A vdd FULL_ADDER_3/XOR_1/w_n16_50# pfet w=16 l=2
+  ad=96 pd=44 as=0 ps=0
M1157 FULL_ADDER_3/XOR_1/a_18_52# FULL_ADDER_3/XOR_1/a_n3_n2# vdd FULL_ADDER_3/XOR_1/w_n16_50# pfet w=16 l=2
+  ad=80 pd=42 as=0 ps=0
M1158 FULL_ADDER_3/SUM FULL_ADDER_3/CIN FULL_ADDER_3/XOR_1/a_18_52# FULL_ADDER_3/XOR_1/w_n16_50# pfet w=16 l=2
+  ad=224 pd=92 as=0 ps=0
M1159 FULL_ADDER_3/XOR_1/a_47_52# FULL_ADDER_3/XOR_1/a_21_19# FULL_ADDER_3/SUM FULL_ADDER_3/XOR_1/w_n16_50# pfet w=16 l=2
+  ad=80 pd=42 as=0 ps=0
M1160 vdd FULL_ADDER_3/XOR_1/a_52_45# FULL_ADDER_3/XOR_1/a_47_52# FULL_ADDER_3/XOR_1/w_n16_50# pfet w=16 l=2
+  ad=0 pd=0 as=0 ps=0
M1161 vdd FULL_ADDER_3/CIN FULL_ADDER_3/XOR_1/a_52_45# FULL_ADDER_3/XOR_1/w_n16_50# pfet w=16 l=2
+  ad=0 pd=0 as=96 ps=44
M1162 FULL_ADDER_3/XOR_1/a_n3_n2# FULL_ADDER_3/XOR_1/A gnd Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1163 FULL_ADDER_3/XOR_1/a_18_n2# FULL_ADDER_3/CIN gnd Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1164 FULL_ADDER_3/SUM FULL_ADDER_3/XOR_1/a_21_19# FULL_ADDER_3/XOR_1/a_18_n2# Gnd nfet w=8 l=2
+  ad=120 pd=62 as=0 ps=0
M1165 FULL_ADDER_3/XOR_1/a_48_n2# FULL_ADDER_3/XOR_1/a_n3_n2# FULL_ADDER_3/SUM Gnd nfet w=8 l=2
+  ad=48 pd=28 as=0 ps=0
M1166 gnd FULL_ADDER_3/XOR_1/a_52_45# FULL_ADDER_3/XOR_1/a_48_n2# Gnd nfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1167 gnd FULL_ADDER_3/CIN FULL_ADDER_3/XOR_1/a_52_45# Gnd nfet w=8 l=2
+  ad=0 pd=0 as=40 ps=26
M1168 FULL_ADDER_3/XOR_0/a_n3_n2# FULL_ADDER_3/XOR_0/A vdd FULL_ADDER_3/XOR_0/w_n16_50# pfet w=16 l=2
+  ad=96 pd=44 as=0 ps=0
M1169 FULL_ADDER_3/XOR_0/a_18_52# FULL_ADDER_3/XOR_0/a_n3_n2# vdd FULL_ADDER_3/XOR_0/w_n16_50# pfet w=16 l=2
+  ad=80 pd=42 as=0 ps=0
M1170 FULL_ADDER_3/XOR_1/A FULL_ADDER_3/B FULL_ADDER_3/XOR_0/a_18_52# FULL_ADDER_3/XOR_0/w_n16_50# pfet w=16 l=2
+  ad=224 pd=92 as=0 ps=0
M1171 FULL_ADDER_3/XOR_0/a_47_52# FULL_ADDER_3/XOR_0/a_21_19# FULL_ADDER_3/XOR_1/A FULL_ADDER_3/XOR_0/w_n16_50# pfet w=16 l=2
+  ad=80 pd=42 as=0 ps=0
M1172 vdd FULL_ADDER_3/XOR_0/a_52_45# FULL_ADDER_3/XOR_0/a_47_52# FULL_ADDER_3/XOR_0/w_n16_50# pfet w=16 l=2
+  ad=0 pd=0 as=0 ps=0
M1173 vdd FULL_ADDER_3/B FULL_ADDER_3/XOR_0/a_52_45# FULL_ADDER_3/XOR_0/w_n16_50# pfet w=16 l=2
+  ad=0 pd=0 as=96 ps=44
M1174 FULL_ADDER_3/XOR_0/a_n3_n2# FULL_ADDER_3/XOR_0/A gnd Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1175 FULL_ADDER_3/XOR_0/a_18_n2# FULL_ADDER_3/B gnd Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1176 FULL_ADDER_3/XOR_1/A FULL_ADDER_3/XOR_0/a_21_19# FULL_ADDER_3/XOR_0/a_18_n2# Gnd nfet w=8 l=2
+  ad=120 pd=62 as=0 ps=0
M1177 FULL_ADDER_3/XOR_0/a_48_n2# FULL_ADDER_3/XOR_0/a_n3_n2# FULL_ADDER_3/XOR_1/A Gnd nfet w=8 l=2
+  ad=48 pd=28 as=0 ps=0
M1178 gnd FULL_ADDER_3/XOR_0/a_52_45# FULL_ADDER_3/XOR_0/a_48_n2# Gnd nfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1179 gnd FULL_ADDER_3/B FULL_ADDER_3/XOR_0/a_52_45# Gnd nfet w=8 l=2
+  ad=0 pd=0 as=40 ps=26
M1180 FULL_ADDER_0/COUT FULL_ADDER_0/NAND_2/IN_A vdd vdd pfet w=16 l=2
+  ad=192 pd=56 as=0 ps=0
M1181 vdd FULL_ADDER_0/NAND_2/IN_B FULL_ADDER_0/COUT vdd pfet w=16 l=2
+  ad=0 pd=0 as=0 ps=0
M1182 FULL_ADDER_0/NAND_2/DS FULL_ADDER_0/NAND_2/IN_A gnd Gnd nfet w=8 l=2
+  ad=96 pd=40 as=0 ps=0
M1183 FULL_ADDER_0/COUT FULL_ADDER_0/NAND_2/IN_B FULL_ADDER_0/NAND_2/DS Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1184 FULL_ADDER_0/NAND_2/IN_B FULL_ADDER_0/B vdd vdd pfet w=16 l=2
+  ad=192 pd=56 as=0 ps=0
M1185 vdd gnd FULL_ADDER_0/NAND_2/IN_B vdd pfet w=16 l=2
+  ad=0 pd=0 as=0 ps=0
M1186 FULL_ADDER_0/NAND_1/DS FULL_ADDER_0/B gnd Gnd nfet w=8 l=2
+  ad=96 pd=40 as=0 ps=0
M1187 FULL_ADDER_0/NAND_2/IN_B gnd FULL_ADDER_0/NAND_1/DS Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1188 FULL_ADDER_0/NAND_2/IN_A FULL_ADDER_0/CIN vdd vdd pfet w=16 l=2
+  ad=192 pd=56 as=0 ps=0
M1189 vdd FULL_ADDER_0/XOR_1/A FULL_ADDER_0/NAND_2/IN_A vdd pfet w=16 l=2
+  ad=0 pd=0 as=0 ps=0
M1190 FULL_ADDER_0/NAND_0/DS FULL_ADDER_0/CIN gnd Gnd nfet w=8 l=2
+  ad=96 pd=40 as=0 ps=0
M1191 FULL_ADDER_0/NAND_2/IN_A FULL_ADDER_0/XOR_1/A FULL_ADDER_0/NAND_0/DS Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1192 FULL_ADDER_0/XOR_1/a_n3_n2# FULL_ADDER_0/XOR_1/A vdd FULL_ADDER_0/XOR_1/w_n16_50# pfet w=16 l=2
+  ad=96 pd=44 as=0 ps=0
M1193 FULL_ADDER_0/XOR_1/a_18_52# FULL_ADDER_0/XOR_1/a_n3_n2# vdd FULL_ADDER_0/XOR_1/w_n16_50# pfet w=16 l=2
+  ad=80 pd=42 as=0 ps=0
M1194 FULL_ADDER_0/SUM FULL_ADDER_0/CIN FULL_ADDER_0/XOR_1/a_18_52# FULL_ADDER_0/XOR_1/w_n16_50# pfet w=16 l=2
+  ad=224 pd=92 as=0 ps=0
M1195 FULL_ADDER_0/XOR_1/a_47_52# FULL_ADDER_0/XOR_1/a_21_19# FULL_ADDER_0/SUM FULL_ADDER_0/XOR_1/w_n16_50# pfet w=16 l=2
+  ad=80 pd=42 as=0 ps=0
M1196 vdd FULL_ADDER_0/XOR_1/a_52_45# FULL_ADDER_0/XOR_1/a_47_52# FULL_ADDER_0/XOR_1/w_n16_50# pfet w=16 l=2
+  ad=0 pd=0 as=0 ps=0
M1197 vdd FULL_ADDER_0/CIN FULL_ADDER_0/XOR_1/a_52_45# FULL_ADDER_0/XOR_1/w_n16_50# pfet w=16 l=2
+  ad=0 pd=0 as=96 ps=44
M1198 FULL_ADDER_0/XOR_1/a_n3_n2# FULL_ADDER_0/XOR_1/A gnd Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1199 FULL_ADDER_0/XOR_1/a_18_n2# FULL_ADDER_0/CIN gnd Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1200 FULL_ADDER_0/SUM FULL_ADDER_0/XOR_1/a_21_19# FULL_ADDER_0/XOR_1/a_18_n2# Gnd nfet w=8 l=2
+  ad=120 pd=62 as=0 ps=0
M1201 FULL_ADDER_0/XOR_1/a_48_n2# FULL_ADDER_0/XOR_1/a_n3_n2# FULL_ADDER_0/SUM Gnd nfet w=8 l=2
+  ad=48 pd=28 as=0 ps=0
M1202 gnd FULL_ADDER_0/XOR_1/a_52_45# FULL_ADDER_0/XOR_1/a_48_n2# Gnd nfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1203 gnd FULL_ADDER_0/CIN FULL_ADDER_0/XOR_1/a_52_45# Gnd nfet w=8 l=2
+  ad=0 pd=0 as=40 ps=26
M1204 FULL_ADDER_0/XOR_0/a_n3_n2# FULL_ADDER_0/XOR_0/A vdd FULL_ADDER_0/XOR_0/w_n16_50# pfet w=16 l=2
+  ad=96 pd=44 as=0 ps=0
M1205 FULL_ADDER_0/XOR_0/a_18_52# FULL_ADDER_0/XOR_0/a_n3_n2# vdd FULL_ADDER_0/XOR_0/w_n16_50# pfet w=16 l=2
+  ad=80 pd=42 as=0 ps=0
M1206 FULL_ADDER_0/XOR_1/A FULL_ADDER_0/B FULL_ADDER_0/XOR_0/a_18_52# FULL_ADDER_0/XOR_0/w_n16_50# pfet w=16 l=2
+  ad=224 pd=92 as=0 ps=0
M1207 FULL_ADDER_0/XOR_0/a_47_52# FULL_ADDER_0/XOR_0/a_21_19# FULL_ADDER_0/XOR_1/A FULL_ADDER_0/XOR_0/w_n16_50# pfet w=16 l=2
+  ad=80 pd=42 as=0 ps=0
M1208 vdd FULL_ADDER_0/XOR_0/a_52_45# FULL_ADDER_0/XOR_0/a_47_52# FULL_ADDER_0/XOR_0/w_n16_50# pfet w=16 l=2
+  ad=0 pd=0 as=0 ps=0
M1209 vdd FULL_ADDER_0/B FULL_ADDER_0/XOR_0/a_52_45# FULL_ADDER_0/XOR_0/w_n16_50# pfet w=16 l=2
+  ad=0 pd=0 as=96 ps=44
M1210 FULL_ADDER_0/XOR_0/a_n3_n2# FULL_ADDER_0/XOR_0/A gnd Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1211 FULL_ADDER_0/XOR_0/a_18_n2# FULL_ADDER_0/B gnd Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1212 FULL_ADDER_0/XOR_1/A FULL_ADDER_0/XOR_0/a_21_19# FULL_ADDER_0/XOR_0/a_18_n2# Gnd nfet w=8 l=2
+  ad=120 pd=62 as=0 ps=0
M1213 FULL_ADDER_0/XOR_0/a_48_n2# FULL_ADDER_0/XOR_0/a_n3_n2# FULL_ADDER_0/XOR_1/A Gnd nfet w=8 l=2
+  ad=48 pd=28 as=0 ps=0
M1214 gnd FULL_ADDER_0/XOR_0/a_52_45# FULL_ADDER_0/XOR_0/a_48_n2# Gnd nfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1215 gnd FULL_ADDER_0/B FULL_ADDER_0/XOR_0/a_52_45# Gnd nfet w=8 l=2
+  ad=0 pd=0 as=40 ps=26
M1216 FULL_ADDER_1/COUT FULL_ADDER_1/NAND_2/IN_A vdd vdd pfet w=16 l=2
+  ad=192 pd=56 as=0 ps=0
M1217 vdd FULL_ADDER_1/NAND_2/IN_B FULL_ADDER_1/COUT vdd pfet w=16 l=2
+  ad=0 pd=0 as=0 ps=0
M1218 FULL_ADDER_1/NAND_2/DS FULL_ADDER_1/NAND_2/IN_A gnd Gnd nfet w=8 l=2
+  ad=96 pd=40 as=0 ps=0
M1219 FULL_ADDER_1/COUT FULL_ADDER_1/NAND_2/IN_B FULL_ADDER_1/NAND_2/DS Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1220 FULL_ADDER_1/NAND_2/IN_B FULL_ADDER_1/B vdd vdd pfet w=16 l=2
+  ad=192 pd=56 as=0 ps=0
M1221 vdd gnd FULL_ADDER_1/NAND_2/IN_B vdd pfet w=16 l=2
+  ad=0 pd=0 as=0 ps=0
M1222 FULL_ADDER_1/NAND_1/DS FULL_ADDER_1/B gnd Gnd nfet w=8 l=2
+  ad=96 pd=40 as=0 ps=0
M1223 FULL_ADDER_1/NAND_2/IN_B gnd FULL_ADDER_1/NAND_1/DS Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1224 FULL_ADDER_1/NAND_2/IN_A FULL_ADDER_1/CIN vdd vdd pfet w=16 l=2
+  ad=192 pd=56 as=0 ps=0
M1225 vdd FULL_ADDER_1/XOR_1/A FULL_ADDER_1/NAND_2/IN_A vdd pfet w=16 l=2
+  ad=0 pd=0 as=0 ps=0
M1226 FULL_ADDER_1/NAND_0/DS FULL_ADDER_1/CIN gnd Gnd nfet w=8 l=2
+  ad=96 pd=40 as=0 ps=0
M1227 FULL_ADDER_1/NAND_2/IN_A FULL_ADDER_1/XOR_1/A FULL_ADDER_1/NAND_0/DS Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1228 FULL_ADDER_1/XOR_1/a_n3_n2# FULL_ADDER_1/XOR_1/A vdd FULL_ADDER_1/XOR_1/w_n16_50# pfet w=16 l=2
+  ad=96 pd=44 as=0 ps=0
M1229 FULL_ADDER_1/XOR_1/a_18_52# FULL_ADDER_1/XOR_1/a_n3_n2# vdd FULL_ADDER_1/XOR_1/w_n16_50# pfet w=16 l=2
+  ad=80 pd=42 as=0 ps=0
M1230 FULL_ADDER_1/SUM FULL_ADDER_1/CIN FULL_ADDER_1/XOR_1/a_18_52# FULL_ADDER_1/XOR_1/w_n16_50# pfet w=16 l=2
+  ad=224 pd=92 as=0 ps=0
M1231 FULL_ADDER_1/XOR_1/a_47_52# FULL_ADDER_1/XOR_1/a_21_19# FULL_ADDER_1/SUM FULL_ADDER_1/XOR_1/w_n16_50# pfet w=16 l=2
+  ad=80 pd=42 as=0 ps=0
M1232 vdd FULL_ADDER_1/XOR_1/a_52_45# FULL_ADDER_1/XOR_1/a_47_52# FULL_ADDER_1/XOR_1/w_n16_50# pfet w=16 l=2
+  ad=0 pd=0 as=0 ps=0
M1233 vdd FULL_ADDER_1/CIN FULL_ADDER_1/XOR_1/a_52_45# FULL_ADDER_1/XOR_1/w_n16_50# pfet w=16 l=2
+  ad=0 pd=0 as=96 ps=44
M1234 FULL_ADDER_1/XOR_1/a_n3_n2# FULL_ADDER_1/XOR_1/A gnd Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1235 FULL_ADDER_1/XOR_1/a_18_n2# FULL_ADDER_1/CIN gnd Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1236 FULL_ADDER_1/SUM FULL_ADDER_1/XOR_1/a_21_19# FULL_ADDER_1/XOR_1/a_18_n2# Gnd nfet w=8 l=2
+  ad=120 pd=62 as=0 ps=0
M1237 FULL_ADDER_1/XOR_1/a_48_n2# FULL_ADDER_1/XOR_1/a_n3_n2# FULL_ADDER_1/SUM Gnd nfet w=8 l=2
+  ad=48 pd=28 as=0 ps=0
M1238 gnd FULL_ADDER_1/XOR_1/a_52_45# FULL_ADDER_1/XOR_1/a_48_n2# Gnd nfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1239 gnd FULL_ADDER_1/CIN FULL_ADDER_1/XOR_1/a_52_45# Gnd nfet w=8 l=2
+  ad=0 pd=0 as=40 ps=26
M1240 FULL_ADDER_1/XOR_0/a_n3_n2# FULL_ADDER_1/XOR_0/A vdd FULL_ADDER_1/XOR_0/w_n16_50# pfet w=16 l=2
+  ad=96 pd=44 as=0 ps=0
M1241 FULL_ADDER_1/XOR_0/a_18_52# FULL_ADDER_1/XOR_0/a_n3_n2# vdd FULL_ADDER_1/XOR_0/w_n16_50# pfet w=16 l=2
+  ad=80 pd=42 as=0 ps=0
M1242 FULL_ADDER_1/XOR_1/A FULL_ADDER_1/B FULL_ADDER_1/XOR_0/a_18_52# FULL_ADDER_1/XOR_0/w_n16_50# pfet w=16 l=2
+  ad=224 pd=92 as=0 ps=0
M1243 FULL_ADDER_1/XOR_0/a_47_52# FULL_ADDER_1/XOR_0/a_21_19# FULL_ADDER_1/XOR_1/A FULL_ADDER_1/XOR_0/w_n16_50# pfet w=16 l=2
+  ad=80 pd=42 as=0 ps=0
M1244 vdd FULL_ADDER_1/XOR_0/a_52_45# FULL_ADDER_1/XOR_0/a_47_52# FULL_ADDER_1/XOR_0/w_n16_50# pfet w=16 l=2
+  ad=0 pd=0 as=0 ps=0
M1245 vdd FULL_ADDER_1/B FULL_ADDER_1/XOR_0/a_52_45# FULL_ADDER_1/XOR_0/w_n16_50# pfet w=16 l=2
+  ad=0 pd=0 as=96 ps=44
M1246 FULL_ADDER_1/XOR_0/a_n3_n2# FULL_ADDER_1/XOR_0/A gnd Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1247 FULL_ADDER_1/XOR_0/a_18_n2# FULL_ADDER_1/B gnd Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1248 FULL_ADDER_1/XOR_1/A FULL_ADDER_1/XOR_0/a_21_19# FULL_ADDER_1/XOR_0/a_18_n2# Gnd nfet w=8 l=2
+  ad=120 pd=62 as=0 ps=0
M1249 FULL_ADDER_1/XOR_0/a_48_n2# FULL_ADDER_1/XOR_0/a_n3_n2# FULL_ADDER_1/XOR_1/A Gnd nfet w=8 l=2
+  ad=48 pd=28 as=0 ps=0
M1250 gnd FULL_ADDER_1/XOR_0/a_52_45# FULL_ADDER_1/XOR_0/a_48_n2# Gnd nfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1251 gnd FULL_ADDER_1/B FULL_ADDER_1/XOR_0/a_52_45# Gnd nfet w=8 l=2
+  ad=0 pd=0 as=40 ps=26
M1252 FULL_ADDER_2/COUT FULL_ADDER_2/NAND_2/IN_A vdd vdd pfet w=16 l=2
+  ad=192 pd=56 as=0 ps=0
M1253 vdd FULL_ADDER_2/NAND_2/IN_B FULL_ADDER_2/COUT vdd pfet w=16 l=2
+  ad=0 pd=0 as=0 ps=0
M1254 FULL_ADDER_2/NAND_2/DS FULL_ADDER_2/NAND_2/IN_A gnd Gnd nfet w=8 l=2
+  ad=96 pd=40 as=0 ps=0
M1255 FULL_ADDER_2/COUT FULL_ADDER_2/NAND_2/IN_B FULL_ADDER_2/NAND_2/DS Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1256 FULL_ADDER_2/NAND_2/IN_B FULL_ADDER_2/B vdd vdd pfet w=16 l=2
+  ad=192 pd=56 as=0 ps=0
M1257 vdd gnd FULL_ADDER_2/NAND_2/IN_B vdd pfet w=16 l=2
+  ad=0 pd=0 as=0 ps=0
M1258 FULL_ADDER_2/NAND_1/DS FULL_ADDER_2/B gnd Gnd nfet w=8 l=2
+  ad=96 pd=40 as=0 ps=0
M1259 FULL_ADDER_2/NAND_2/IN_B gnd FULL_ADDER_2/NAND_1/DS Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1260 FULL_ADDER_2/NAND_2/IN_A FULL_ADDER_2/CIN vdd vdd pfet w=16 l=2
+  ad=192 pd=56 as=0 ps=0
M1261 vdd FULL_ADDER_2/XOR_1/A FULL_ADDER_2/NAND_2/IN_A vdd pfet w=16 l=2
+  ad=0 pd=0 as=0 ps=0
M1262 FULL_ADDER_2/NAND_0/DS FULL_ADDER_2/CIN gnd Gnd nfet w=8 l=2
+  ad=96 pd=40 as=0 ps=0
M1263 FULL_ADDER_2/NAND_2/IN_A FULL_ADDER_2/XOR_1/A FULL_ADDER_2/NAND_0/DS Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1264 FULL_ADDER_2/XOR_1/a_n3_n2# FULL_ADDER_2/XOR_1/A vdd FULL_ADDER_2/XOR_1/w_n16_50# pfet w=16 l=2
+  ad=96 pd=44 as=0 ps=0
M1265 FULL_ADDER_2/XOR_1/a_18_52# FULL_ADDER_2/XOR_1/a_n3_n2# vdd FULL_ADDER_2/XOR_1/w_n16_50# pfet w=16 l=2
+  ad=80 pd=42 as=0 ps=0
M1266 FULL_ADDER_2/SUM FULL_ADDER_2/CIN FULL_ADDER_2/XOR_1/a_18_52# FULL_ADDER_2/XOR_1/w_n16_50# pfet w=16 l=2
+  ad=224 pd=92 as=0 ps=0
M1267 FULL_ADDER_2/XOR_1/a_47_52# FULL_ADDER_2/XOR_1/a_21_19# FULL_ADDER_2/SUM FULL_ADDER_2/XOR_1/w_n16_50# pfet w=16 l=2
+  ad=80 pd=42 as=0 ps=0
M1268 vdd FULL_ADDER_2/XOR_1/a_52_45# FULL_ADDER_2/XOR_1/a_47_52# FULL_ADDER_2/XOR_1/w_n16_50# pfet w=16 l=2
+  ad=0 pd=0 as=0 ps=0
M1269 vdd FULL_ADDER_2/CIN FULL_ADDER_2/XOR_1/a_52_45# FULL_ADDER_2/XOR_1/w_n16_50# pfet w=16 l=2
+  ad=0 pd=0 as=96 ps=44
M1270 FULL_ADDER_2/XOR_1/a_n3_n2# FULL_ADDER_2/XOR_1/A gnd Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1271 FULL_ADDER_2/XOR_1/a_18_n2# FULL_ADDER_2/CIN gnd Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1272 FULL_ADDER_2/SUM FULL_ADDER_2/XOR_1/a_21_19# FULL_ADDER_2/XOR_1/a_18_n2# Gnd nfet w=8 l=2
+  ad=120 pd=62 as=0 ps=0
M1273 FULL_ADDER_2/XOR_1/a_48_n2# FULL_ADDER_2/XOR_1/a_n3_n2# FULL_ADDER_2/SUM Gnd nfet w=8 l=2
+  ad=48 pd=28 as=0 ps=0
M1274 gnd FULL_ADDER_2/XOR_1/a_52_45# FULL_ADDER_2/XOR_1/a_48_n2# Gnd nfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1275 gnd FULL_ADDER_2/CIN FULL_ADDER_2/XOR_1/a_52_45# Gnd nfet w=8 l=2
+  ad=0 pd=0 as=40 ps=26
M1276 FULL_ADDER_2/XOR_0/a_n3_n2# FULL_ADDER_2/XOR_0/A vdd FULL_ADDER_2/XOR_0/w_n16_50# pfet w=16 l=2
+  ad=96 pd=44 as=0 ps=0
M1277 FULL_ADDER_2/XOR_0/a_18_52# FULL_ADDER_2/XOR_0/a_n3_n2# vdd FULL_ADDER_2/XOR_0/w_n16_50# pfet w=16 l=2
+  ad=80 pd=42 as=0 ps=0
M1278 FULL_ADDER_2/XOR_1/A FULL_ADDER_2/B FULL_ADDER_2/XOR_0/a_18_52# FULL_ADDER_2/XOR_0/w_n16_50# pfet w=16 l=2
+  ad=224 pd=92 as=0 ps=0
M1279 FULL_ADDER_2/XOR_0/a_47_52# FULL_ADDER_2/XOR_0/a_21_19# FULL_ADDER_2/XOR_1/A FULL_ADDER_2/XOR_0/w_n16_50# pfet w=16 l=2
+  ad=80 pd=42 as=0 ps=0
M1280 vdd FULL_ADDER_2/XOR_0/a_52_45# FULL_ADDER_2/XOR_0/a_47_52# FULL_ADDER_2/XOR_0/w_n16_50# pfet w=16 l=2
+  ad=0 pd=0 as=0 ps=0
M1281 vdd FULL_ADDER_2/B FULL_ADDER_2/XOR_0/a_52_45# FULL_ADDER_2/XOR_0/w_n16_50# pfet w=16 l=2
+  ad=0 pd=0 as=96 ps=44
M1282 FULL_ADDER_2/XOR_0/a_n3_n2# FULL_ADDER_2/XOR_0/A gnd Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1283 FULL_ADDER_2/XOR_0/a_18_n2# FULL_ADDER_2/B gnd Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1284 FULL_ADDER_2/XOR_1/A FULL_ADDER_2/XOR_0/a_21_19# FULL_ADDER_2/XOR_0/a_18_n2# Gnd nfet w=8 l=2
+  ad=120 pd=62 as=0 ps=0
M1285 FULL_ADDER_2/XOR_0/a_48_n2# FULL_ADDER_2/XOR_0/a_n3_n2# FULL_ADDER_2/XOR_1/A Gnd nfet w=8 l=2
+  ad=48 pd=28 as=0 ps=0
M1286 gnd FULL_ADDER_2/XOR_0/a_52_45# FULL_ADDER_2/XOR_0/a_48_n2# Gnd nfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1287 gnd FULL_ADDER_2/B FULL_ADDER_2/XOR_0/a_52_45# Gnd nfet w=8 l=2
+  ad=0 pd=0 as=40 ps=26
C0 vdd FULL_ADDER_0/NAND_2/IN_B 8.5fF
C1 vdd FULL_ADDER_5/NAND_2/IN_A 25.0fF
C2 vdd FULL_ADDER_2/XOR_1/A 4.6fF
C3 vdd FULL_ADDER_0/XOR_1/A 4.6fF
C4 vdd FULL_ADDER_0/NAND_2/IN_A 25.0fF
C5 FULL_ADDER_1/XOR_0/w_n16_50# FULL_ADDER_1/B 4.4fF
C6 FULL_ADDER_3/XOR_0/w_n16_50# FULL_ADDER_3/B 4.4fF
C7 vdd FULL_ADDER_4/XOR_1/w_n16_50# 8.5fF
C8 vdd FULL_ADDER_5/NAND_2/IN_B 8.5fF
C9 FULL_ADDER_7/XOR_1/A vdd 4.6fF
C10 vdd FULL_ADDER_2/XOR_0/w_n16_50# 16.4fF
C11 vdd FULL_ADDER_0/XOR_0/w_n16_50# 16.4fF
C12 vdd FULL_ADDER_3/NAND_2/IN_B 8.5fF
C13 vdd FULL_ADDER_4/NAND_2/IN_A 25.0fF
C14 vdd FULL_ADDER_1/CIN 11.8fF
C15 vdd FULL_ADDER_1/XOR_1/A 4.6fF
C16 vdd FULL_ADDER_7/XOR_0/w_n16_50# 16.4fF
C17 vdd FULL_ADDER_4/CIN 11.8fF
C18 vdd FULL_ADDER_2/B 8.5fF
C19 vdd FULL_ADDER_6/NAND_2/IN_B 8.5fF
C20 vdd FULL_ADDER_0/B 8.5fF
C21 FULL_ADDER_3/XOR_1/w_n16_50# FULL_ADDER_3/CIN 4.4fF
C22 FULL_ADDER_5/XOR_0/w_n16_50# FULL_ADDER_5/B 4.4fF
C23 FULL_ADDER_7/NAND_2/IN_B vdd 8.5fF
C24 vdd FULL_ADDER_7/B 8.5fF
C25 vdd FULL_ADDER_1/NAND_2/IN_A 25.0fF
C26 vdd FULL_ADDER_6/B 8.5fF
C27 FULL_ADDER_7/NAND_2/IN_A vdd 25.0fF
C28 vdd FULL_ADDER_3/XOR_1/w_n16_50# 8.5fF
C29 vdd FULL_ADDER_5/XOR_0/w_n16_50# 16.4fF
C30 FULL_ADDER_1/XOR_1/w_n16_50# FULL_ADDER_1/CIN 4.4fF
C31 FULL_ADDER_6/XOR_1/w_n16_50# FULL_ADDER_6/CIN 4.4fF
C32 vdd FULL_ADDER_4/XOR_1/A 4.6fF
C33 vdd FULL_ADDER_6/XOR_1/w_n16_50# 8.5fF
C34 vdd FULL_ADDER_5/XOR_1/w_n16_50# 8.5fF
C35 FULL_ADDER_5/XOR_1/w_n16_50# FULL_ADDER_5/CIN 4.4fF
C36 vdd FULL_ADDER_0/XOR_1/w_n16_50# 8.5fF
C37 FULL_ADDER_6/XOR_0/w_n16_50# FULL_ADDER_6/B 4.4fF
C38 vdd FULL_ADDER_4/XOR_0/w_n16_50# 16.4fF
C39 vdd FULL_ADDER_4/NAND_2/IN_B 8.5fF
C40 vdd FULL_ADDER_2/NAND_2/IN_B 8.5fF
C41 FULL_ADDER_0/XOR_1/w_n16_50# FULL_ADDER_0/CIN 4.4fF
C42 FULL_ADDER_4/XOR_0/w_n16_50# FULL_ADDER_4/B 4.4fF
C43 vdd FULL_ADDER_3/CIN 11.8fF
C44 vdd FULL_ADDER_5/B 8.5fF
C45 vdd FULL_ADDER_2/XOR_1/w_n16_50# 8.5fF
C46 FULL_ADDER_4/XOR_1/w_n16_50# FULL_ADDER_4/CIN 4.4fF
C47 vdd FULL_ADDER_6/CIN 11.8fF
C48 FULL_ADDER_7/XOR_1/w_n16_50# vdd 8.5fF
C49 vdd FULL_ADDER_3/XOR_1/A 4.6fF
C50 vdd FULL_ADDER_5/CIN 11.8fF
C51 FULL_ADDER_2/XOR_0/w_n16_50# FULL_ADDER_2/B 4.4fF
C52 FULL_ADDER_0/XOR_0/w_n16_50# FULL_ADDER_0/B 4.4fF
C53 vdd FULL_ADDER_0/CIN 11.8fF
C54 vdd FULL_ADDER_4/B 8.5fF
C55 vdd FULL_ADDER_1/XOR_0/w_n16_50# 16.4fF
C56 vdd FULL_ADDER_3/XOR_0/w_n16_50# 16.4fF
C57 vdd FULL_ADDER_6/XOR_1/A 4.6fF
C58 FULL_ADDER_2/XOR_1/w_n16_50# FULL_ADDER_2/CIN 4.4fF
C59 vdd FULL_ADDER_1/NAND_2/IN_B 8.5fF
C60 vdd FULL_ADDER_2/NAND_2/IN_A 25.0fF
C61 FULL_ADDER_7/CIN vdd 11.8fF
C62 FULL_ADDER_7/XOR_1/w_n16_50# FULL_ADDER_7/CIN 4.4fF
C63 vdd FULL_ADDER_3/NAND_2/IN_A 25.0fF
C64 vdd FULL_ADDER_2/CIN 11.8fF
C65 vdd FULL_ADDER_6/XOR_0/w_n16_50# 16.4fF
C66 vdd FULL_ADDER_6/NAND_2/IN_A 25.0fF
C67 vdd FULL_ADDER_5/XOR_1/A 4.6fF
C68 FULL_ADDER_7/XOR_0/w_n16_50# FULL_ADDER_7/B 4.4fF
C69 vdd FULL_ADDER_1/XOR_1/w_n16_50# 8.5fF
C70 vdd FULL_ADDER_1/B 8.5fF
C71 vdd FULL_ADDER_3/B 8.5fF
C72 FULL_ADDER_2/m2_n16_58# gnd! 3.8fF **FLOATING
C73 FULL_ADDER_2/A gnd! 10.1fF **FLOATING
C74 FULL_ADDER_2/XOR_0/a_52_45# gnd! 21.0fF
C75 FULL_ADDER_2/XOR_0/a_21_19# gnd! 19.0fF
C76 FULL_ADDER_2/XOR_0/a_n3_n2# gnd! 38.4fF
C77 FULL_ADDER_2/XOR_0/A gnd! 26.0fF
C78 FULL_ADDER_2/B gnd! 243.4fF
C79 FULL_ADDER_2/SUM gnd! 26.4fF
C80 FULL_ADDER_2/XOR_1/a_52_45# gnd! 21.0fF
C81 FULL_ADDER_2/XOR_1/a_21_19# gnd! 19.0fF
C82 FULL_ADDER_2/XOR_1/a_n3_n2# gnd! 38.4fF
C83 FULL_ADDER_2/XOR_1/A gnd! 71.5fF
C84 FULL_ADDER_2/CIN gnd! 101.1fF
C85 FULL_ADDER_2/NAND_2/IN_A gnd! 21.4fF
C86 FULL_ADDER_2/COUT gnd! 37.9fF
C87 FULL_ADDER_2/NAND_2/IN_B gnd! 30.0fF
C88 FULL_ADDER_1/m2_n16_58# gnd! 3.8fF **FLOATING
C89 FULL_ADDER_1/A gnd! 10.1fF **FLOATING
C90 FULL_ADDER_1/XOR_0/a_52_45# gnd! 21.0fF
C91 FULL_ADDER_1/XOR_0/a_21_19# gnd! 19.0fF
C92 FULL_ADDER_1/XOR_0/a_n3_n2# gnd! 38.4fF
C93 FULL_ADDER_1/XOR_0/A gnd! 26.0fF
C94 FULL_ADDER_1/B gnd! 243.4fF
C95 FULL_ADDER_1/SUM gnd! 26.4fF
C96 FULL_ADDER_1/XOR_1/a_52_45# gnd! 21.0fF
C97 FULL_ADDER_1/XOR_1/a_21_19# gnd! 19.0fF
C98 FULL_ADDER_1/XOR_1/a_n3_n2# gnd! 38.4fF
C99 FULL_ADDER_1/XOR_1/A gnd! 71.5fF
C100 FULL_ADDER_1/CIN gnd! 101.1fF
C101 FULL_ADDER_1/NAND_2/IN_A gnd! 21.4fF
C102 FULL_ADDER_1/COUT gnd! 37.9fF
C103 FULL_ADDER_1/NAND_2/IN_B gnd! 30.0fF
C104 FULL_ADDER_0/m2_n16_58# gnd! 3.8fF **FLOATING
C105 FULL_ADDER_0/A gnd! 10.1fF **FLOATING
C106 FULL_ADDER_0/XOR_0/a_52_45# gnd! 21.0fF
C107 FULL_ADDER_0/XOR_0/a_21_19# gnd! 19.0fF
C108 FULL_ADDER_0/XOR_0/a_n3_n2# gnd! 38.4fF
C109 FULL_ADDER_0/XOR_0/A gnd! 26.0fF
C110 FULL_ADDER_0/B gnd! 243.4fF
C111 FULL_ADDER_0/SUM gnd! 26.4fF
C112 FULL_ADDER_0/XOR_1/a_52_45# gnd! 21.0fF
C113 FULL_ADDER_0/XOR_1/a_21_19# gnd! 19.0fF
C114 FULL_ADDER_0/XOR_1/a_n3_n2# gnd! 38.4fF
C115 FULL_ADDER_0/XOR_1/A gnd! 71.5fF
C116 FULL_ADDER_0/CIN gnd! 101.1fF
C117 FULL_ADDER_0/NAND_2/IN_A gnd! 21.4fF
C118 FULL_ADDER_0/COUT gnd! 37.9fF
C119 FULL_ADDER_0/NAND_2/IN_B gnd! 30.0fF
C120 FULL_ADDER_3/m2_n16_58# gnd! 3.8fF **FLOATING
C121 FULL_ADDER_3/A gnd! 10.1fF **FLOATING
C122 FULL_ADDER_3/XOR_0/a_52_45# gnd! 21.0fF
C123 FULL_ADDER_3/XOR_0/a_21_19# gnd! 19.0fF
C124 FULL_ADDER_3/XOR_0/a_n3_n2# gnd! 38.4fF
C125 FULL_ADDER_3/XOR_0/A gnd! 26.0fF
C126 FULL_ADDER_3/B gnd! 243.4fF
C127 FULL_ADDER_3/SUM gnd! 26.4fF
C128 FULL_ADDER_3/XOR_1/a_52_45# gnd! 21.0fF
C129 FULL_ADDER_3/XOR_1/a_21_19# gnd! 19.0fF
C130 FULL_ADDER_3/XOR_1/a_n3_n2# gnd! 38.4fF
C131 FULL_ADDER_3/XOR_1/A gnd! 71.5fF
C132 FULL_ADDER_3/CIN gnd! 101.1fF
C133 FULL_ADDER_3/NAND_2/IN_A gnd! 21.4fF
C134 FULL_ADDER_3/COUT gnd! 37.9fF
C135 FULL_ADDER_3/NAND_2/IN_B gnd! 30.0fF
C136 FULL_ADDER_4/m2_n16_58# gnd! 3.8fF **FLOATING
C137 FULL_ADDER_4/A gnd! 10.1fF **FLOATING
C138 FULL_ADDER_4/XOR_0/a_52_45# gnd! 21.0fF
C139 FULL_ADDER_4/XOR_0/a_21_19# gnd! 19.0fF
C140 FULL_ADDER_4/XOR_0/a_n3_n2# gnd! 38.4fF
C141 FULL_ADDER_4/XOR_0/A gnd! 26.0fF
C142 FULL_ADDER_4/B gnd! 243.4fF
C143 FULL_ADDER_4/SUM gnd! 26.4fF
C144 FULL_ADDER_4/XOR_1/a_52_45# gnd! 21.0fF
C145 FULL_ADDER_4/XOR_1/a_21_19# gnd! 19.0fF
C146 FULL_ADDER_4/XOR_1/a_n3_n2# gnd! 38.4fF
C147 FULL_ADDER_4/XOR_1/A gnd! 71.5fF
C148 FULL_ADDER_4/CIN gnd! 101.1fF
C149 FULL_ADDER_4/NAND_2/IN_A gnd! 21.4fF
C150 FULL_ADDER_4/COUT gnd! 37.9fF
C151 FULL_ADDER_4/NAND_2/IN_B gnd! 30.0fF
C152 FULL_ADDER_5/m2_n16_58# gnd! 3.8fF **FLOATING
C153 FULL_ADDER_5/A gnd! 10.1fF **FLOATING
C154 FULL_ADDER_5/XOR_0/a_52_45# gnd! 21.0fF
C155 FULL_ADDER_5/XOR_0/a_21_19# gnd! 19.0fF
C156 FULL_ADDER_5/XOR_0/a_n3_n2# gnd! 38.4fF
C157 FULL_ADDER_5/XOR_0/A gnd! 26.0fF
C158 FULL_ADDER_5/B gnd! 243.4fF
C159 FULL_ADDER_5/SUM gnd! 26.4fF
C160 FULL_ADDER_5/XOR_1/a_52_45# gnd! 21.0fF
C161 FULL_ADDER_5/XOR_1/a_21_19# gnd! 19.0fF
C162 FULL_ADDER_5/XOR_1/a_n3_n2# gnd! 38.4fF
C163 FULL_ADDER_5/XOR_1/A gnd! 71.5fF
C164 FULL_ADDER_5/CIN gnd! 101.1fF
C165 FULL_ADDER_5/NAND_2/IN_A gnd! 21.4fF
C166 FULL_ADDER_5/COUT gnd! 37.9fF
C167 FULL_ADDER_5/NAND_2/IN_B gnd! 30.0fF
C168 FULL_ADDER_6/m2_n16_58# gnd! 3.8fF **FLOATING
C169 FULL_ADDER_6/A gnd! 10.1fF **FLOATING
C170 FULL_ADDER_6/XOR_0/a_52_45# gnd! 21.0fF
C171 FULL_ADDER_6/XOR_0/a_21_19# gnd! 19.0fF
C172 FULL_ADDER_6/XOR_0/a_n3_n2# gnd! 38.4fF
C173 FULL_ADDER_6/XOR_0/A gnd! 26.0fF
C174 FULL_ADDER_6/B gnd! 243.4fF
C175 FULL_ADDER_6/SUM gnd! 26.4fF
C176 FULL_ADDER_6/XOR_1/a_52_45# gnd! 21.0fF
C177 FULL_ADDER_6/XOR_1/a_21_19# gnd! 19.0fF
C178 FULL_ADDER_6/XOR_1/a_n3_n2# gnd! 38.4fF
C179 FULL_ADDER_6/XOR_1/A gnd! 71.5fF
C180 FULL_ADDER_6/CIN gnd! 101.1fF
C181 FULL_ADDER_6/NAND_2/IN_A gnd! 21.4fF
C182 FULL_ADDER_6/COUT gnd! 37.9fF
C183 FULL_ADDER_6/NAND_2/IN_B gnd! 30.0fF
C184 FULL_ADDER_7/m2_n16_58# gnd! 3.8fF **FLOATING
C185 FULL_ADDER_7/A gnd! 10.1fF **FLOATING
C186 FULL_ADDER_7/XOR_0/a_52_45# gnd! 21.0fF
C187 FULL_ADDER_7/XOR_0/a_21_19# gnd! 19.0fF
C188 FULL_ADDER_7/XOR_0/a_n3_n2# gnd! 38.4fF
C189 FULL_ADDER_7/XOR_0/A gnd! 26.0fF
C190 FULL_ADDER_7/B gnd! 243.4fF
C191 FULL_ADDER_7/SUM gnd! 26.4fF
C192 vdd gnd! 3956.8fF
C193 FULL_ADDER_7/XOR_1/a_52_45# gnd! 21.0fF
C194 FULL_ADDER_7/XOR_1/a_21_19# gnd! 19.0fF
C195 FULL_ADDER_7/XOR_1/a_n3_n2# gnd! 38.4fF
C196 FULL_ADDER_7/XOR_1/A gnd! 71.5fF
C197 FULL_ADDER_7/CIN gnd! 101.1fF
C198 FULL_ADDER_7/NAND_2/IN_A gnd! 21.4fF
C199 FULL_ADDER_7/COUT gnd! 37.9fF
C200 FULL_ADDER_7/NAND_2/IN_B gnd! 30.0fF
