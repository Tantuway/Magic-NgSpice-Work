magic
tech scmos
timestamp 1569418921
<< metal1 >>
rect -60 60 49 67
rect -60 41 -12 60
rect -60 15 -36 41
rect -17 30 -16 34
rect -23 24 -17 27
rect -19 23 -17 24
rect 15 26 23 27
rect 20 23 23 26
rect -114 -5 -36 15
rect -15 7 49 8
rect -114 -77 -90 -5
rect -79 -13 -67 -8
rect -60 -18 -36 -5
rect -32 -6 49 7
rect -32 -65 -24 -6
rect 8 -31 24 -27
rect 19 -38 22 -34
rect 60 -38 78 -34
rect -38 -74 -24 -65
rect -15 -71 49 -65
rect -14 -77 10 -71
rect -114 -92 10 -77
<< metal2 >>
rect -134 30 -21 34
rect 12 30 18 34
rect 46 30 93 34
rect -134 -12 -83 -8
rect -86 -13 -83 -12
rect -75 -45 -71 30
rect -23 24 -19 25
rect -23 -8 -19 20
rect 15 -1 20 22
rect 15 -5 55 -1
rect -63 -13 -19 -8
rect -23 -28 -19 -13
rect -23 -32 -17 -28
rect 51 -34 55 -5
rect 59 -20 63 30
rect 59 -25 74 -20
rect -23 -40 -19 -36
rect 50 -38 56 -34
rect -75 -49 -63 -45
rect -23 -46 -18 -40
rect -36 -50 -18 -46
rect -53 -70 -41 -69
rect -53 -74 -49 -70
rect -45 -74 -41 -70
rect -53 -106 -41 -74
rect 15 -76 19 -38
rect 69 -76 74 -25
rect 82 -38 93 -34
rect 15 -80 74 -76
<< m2contact >>
rect -21 30 -17 34
rect 8 30 12 34
rect 18 30 22 34
rect -23 20 -19 24
rect 15 22 20 26
rect -83 -13 -79 -8
rect -67 -13 -63 -8
rect -63 -49 -59 -45
rect -40 -50 -36 -46
rect -17 -32 -13 -28
rect -19 -40 -15 -36
rect 15 -38 19 -34
rect 46 -38 50 -34
rect 56 -38 60 -34
rect 78 -38 82 -34
rect -49 -74 -45 -70
use NAND  NAND_0
timestamp 1569392509
transform 1 0 -9 0 1 34
box -8 -34 21 34
use NAND  NAND_1
timestamp 1569392509
transform 1 0 29 0 1 34
box -8 -34 21 34
use Inverter  Inverter_0
timestamp 1569345144
transform 1 0 -56 0 1 -43
box -4 -31 20 31
use NAND  NAND_2
timestamp 1569392509
transform 1 0 -9 0 -1 -39
box -8 -34 21 34
use NAND  NAND_3
timestamp 1569392509
transform 1 0 29 0 -1 -38
box -8 -34 21 34
<< labels >>
rlabel metal2 -134 30 -134 34 3 D
rlabel metal2 -134 -12 -134 -8 3 CLK
rlabel metal2 93 30 93 34 7 Q
rlabel metal2 93 -38 93 -34 7 QBAR
rlabel metal2 -53 -106 -41 -106 1 gnd!
<< end >>
