magic
tech scmos
timestamp 1569387030
<< polysilicon >>
rect -49 39 -41 43
rect -37 39 54 43
rect 52 35 54 39
rect -41 33 54 35
rect -41 31 -39 33
rect -41 29 54 31
rect 52 27 54 29
rect -41 25 54 27
rect -41 23 -39 25
rect -41 21 54 23
rect 52 19 54 21
rect -41 17 54 19
rect -41 15 -39 17
rect -41 13 54 15
rect 52 11 54 13
rect -41 9 54 11
rect -41 7 -39 9
rect -41 5 54 7
rect 52 3 54 5
rect -41 1 54 3
rect -41 -1 -39 1
rect -41 -3 54 -1
rect 52 -5 54 -3
rect -41 -7 54 -5
rect -41 -9 -39 -7
rect -41 -11 54 -9
rect 52 -13 54 -11
rect -41 -15 54 -13
rect -41 -17 -39 -15
rect -41 -19 54 -17
rect 52 -23 54 -19
rect -49 -27 -41 -23
rect -37 -27 54 -23
<< metal1 >>
rect -49 39 -41 43
rect -49 -27 -41 -23
<< polycontact >>
rect -41 39 -37 43
rect -41 -27 -37 -23
<< glass >>
rect -52 -31 63 45
<< labels >>
rlabel metal1 -49 39 -49 43 4 a
rlabel metal1 -49 -27 -49 -23 2 b
<< end >>
